** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/OP_AMP_SKY130NM/OP_AMP.sch
**.subckt OP_AMP VSS VDD_1V8 VIN VIP VO LPO LPI
*.ipin VSS
*.ipin VDD_1V8
*.ipin VIN
*.ipin VIP
*.opin VO
*.opin LPO
*.ipin LPI
x1 P5 P2 VSS VSS CNRATR_NCH_4C2F0
x2 P2 P2 VSS VSS CNRATR_NCH_2C8F0
x3 P5 VIN V_TAIL V_TAIL CNRATR_PCH_4C4F0
x4 P2 VIP V_TAIL V_TAIL CNRATR_PCH_4C4F0
x5 V_TAIL P3 VDD_1V8 VDD_1V8 CNRATR_PCH_4C4F0
x6 LPO P3 VDD_1V8 net1 CNRATR_PCH_4C4F0
x7 LPO P2 VSS net2 CNRATR_NCH_4C2F0
x8 P4 P3 VDD_1V8 VDD_1V8 CNRATR_PCH_4C4F0
R1 P4 VSS 2k m=1
XC1 VO VSS sky130_fd_pr__cap_mim_m3_1 W=10 L=100 MF=1 m=1
**.ends

* expanding   symbol:  CNR_ATR_SKY130NM/CNRATR_NCH_4C2F0.sym # of pins=4
** sym_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_4C2F0.sym
** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_4C2F0.sch
.subckt CNRATR_NCH_4C2F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.54 W=3.84 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  CNR_ATR_SKY130NM/CNRATR_NCH_2C8F0.sym # of pins=4
** sym_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_2C8F0.sym
** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_2C8F0.sch
.subckt CNRATR_NCH_2C8F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=2.7 W=1.92 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  CNR_ATR_SKY130NM/CNRATR_PCH_4C4F0.sym # of pins=4
** sym_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_4C4F0.sym
** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_4C4F0.sch
.subckt CNRATR_PCH_4C4F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=1.26 W=3.84 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end

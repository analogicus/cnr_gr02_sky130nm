.param mc_mm_switch=0
.param mc_pr_switch=0

.include tt.spi
.lib "../../../tech/ngspice/temperature.spi" Tl
.lib "../../../tech/ngspice/supply.spi" Vl

.option savecurrents
.save all
.control

optran 0 0 0 10n 10u 0
op
write TB_OTA.raw
exit
.endc
.end

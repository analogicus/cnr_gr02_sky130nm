magic
tech sky130B
magscale 1 2
timestamp 1713553704
<< nwell >>
rect 249 2698 5025 2704
rect 249 1626 5026 2698
<< locali >>
rect 1915 2784 7213 2830
rect 2052 2572 2086 2784
rect 2527 2529 2573 2784
rect 3114 2572 3148 2784
rect 1924 2426 2062 2504
rect 3142 2420 3330 2538
rect 3843 2533 3889 2784
rect 4384 2568 4418 2784
rect 2512 1934 2606 2390
rect 3114 2179 3148 2364
rect 3114 2145 3223 2179
rect 3189 1963 3223 2145
rect 3756 1928 3940 2390
rect 4384 2239 4418 2360
rect 4384 2205 4619 2239
rect 4585 1951 4619 2205
rect 1822 1834 1960 1912
rect 3220 1800 3334 1892
rect 2426 1469 2500 1799
rect 2426 1407 2432 1469
rect 2494 1407 2500 1469
rect 2426 1401 2500 1407
rect 2192 1124 2570 1248
rect 1828 540 1972 806
rect 2872 518 3016 784
rect 2242 96 2750 240
rect 0 20 96 96
rect 1734 20 7742 96
rect 0 -158 7742 20
rect 462 -304 810 -180
rect 1780 -294 2128 -170
rect 3084 -304 3432 -180
rect 4362 -294 4710 -170
rect 5598 -308 5946 -184
rect 6940 -304 7288 -180
rect 7646 -264 7742 -158
rect 462 -1328 810 -1204
rect 1758 -1320 2106 -1196
rect 3058 -1320 3406 -1196
rect 4358 -1310 4706 -1186
rect 5620 -1320 5968 -1196
rect 6948 -1314 7296 -1190
<< viali >>
rect 641 1577 683 1619
rect 2432 1407 2494 1469
<< metal1 >>
rect 3003 2266 3055 2444
rect 1814 2214 3055 2266
rect 3081 1625 3135 1840
rect 629 1619 3135 1625
rect 629 1577 641 1619
rect 683 1577 3135 1619
rect 629 1571 3135 1577
rect 2426 1469 2500 1481
rect 2426 1407 2432 1469
rect 2494 1407 2500 1469
rect 2426 976 2500 1407
rect 2408 906 2500 976
rect 2426 879 2500 906
rect 654 -976 6834 -546
use M9  M9_0
timestamp 1713524830
transform 0 1 2600 -1 0 2468
box -236 -584 236 584
use M9  M9_1
timestamp 1713524830
transform 0 1 3870 -1 0 2464
box -236 -584 236 584
use M10  M10_0
timestamp 1713518505
transform 0 1 2580 -1 0 1864
box -236 -684 236 684
use M10  M10_1
timestamp 1713518505
transform 0 1 3970 -1 0 1860
box -236 -684 236 684
use p4  p4_0
timestamp 1713553704
transform 1 0 0 0 1 0
box 0 0 1980 2830
use Q1  Q1_0 ../design/CNR_GR02_SKY130NM
timestamp 1713553704
transform 1 0 -12 0 1 -2016
box 0 600 7780 1940
use Q2  Q2_0
timestamp 1713553704
transform 1 0 -6028 0 1 -586
box 7780 600 9120 1940
<< end >>

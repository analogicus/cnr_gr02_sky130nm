magic
tech sky130B
magscale 1 2
timestamp 1713258222
<< error_p >>
rect -88 231 -30 237
rect 30 231 88 237
rect -88 197 -76 231
rect 30 197 42 231
rect -88 191 -30 197
rect 30 191 88 197
rect -88 -197 -30 -191
rect 30 -197 88 -191
rect -88 -231 -76 -197
rect 30 -231 42 -197
rect -88 -237 -30 -231
rect 30 -237 88 -231
<< nwell >>
rect -285 -369 285 369
<< pmos >>
rect -89 -150 -29 150
rect 29 -150 89 150
<< pdiff >>
rect -147 138 -89 150
rect -147 -138 -135 138
rect -101 -138 -89 138
rect -147 -150 -89 -138
rect -29 138 29 150
rect -29 -138 -17 138
rect 17 -138 29 138
rect -29 -150 29 -138
rect 89 138 147 150
rect 89 -138 101 138
rect 135 -138 147 138
rect 89 -150 147 -138
<< pdiffc >>
rect -135 -138 -101 138
rect -17 -138 17 138
rect 101 -138 135 138
<< nsubdiff >>
rect -249 299 -153 333
rect 153 299 249 333
rect -249 237 -215 299
rect 215 237 249 299
rect -249 -299 -215 -237
rect 215 -299 249 -237
rect -249 -333 -153 -299
rect 153 -333 249 -299
<< nsubdiffcont >>
rect -153 299 153 333
rect -249 -237 -215 237
rect 215 -237 249 237
rect -153 -333 153 -299
<< poly >>
rect -92 231 -26 247
rect -92 197 -76 231
rect -42 197 -26 231
rect -92 181 -26 197
rect 26 231 92 247
rect 26 197 42 231
rect 76 197 92 231
rect 26 181 92 197
rect -89 150 -29 181
rect 29 150 89 181
rect -89 -181 -29 -150
rect 29 -181 89 -150
rect -92 -197 -26 -181
rect -92 -231 -76 -197
rect -42 -231 -26 -197
rect -92 -247 -26 -231
rect 26 -197 92 -181
rect 26 -231 42 -197
rect 76 -231 92 -197
rect 26 -247 92 -231
<< polycont >>
rect -76 197 -42 231
rect 42 197 76 231
rect -76 -231 -42 -197
rect 42 -231 76 -197
<< locali >>
rect -249 299 -153 333
rect 153 299 249 333
rect -249 237 -215 299
rect 215 237 249 299
rect -92 197 -76 231
rect -42 197 -26 231
rect 26 197 42 231
rect 76 197 92 231
rect -135 138 -101 154
rect -135 -154 -101 -138
rect -17 138 17 154
rect -17 -154 17 -138
rect 101 138 135 154
rect 101 -154 135 -138
rect -92 -231 -76 -197
rect -42 -231 -26 -197
rect 26 -231 42 -197
rect 76 -231 92 -197
rect -249 -299 -215 -237
rect 215 -299 249 -237
rect -249 -333 -153 -299
rect 153 -333 249 -299
<< viali >>
rect -76 197 -42 231
rect 42 197 76 231
rect -135 -138 -101 138
rect -17 -138 17 138
rect 101 -138 135 138
rect -76 -231 -42 -197
rect 42 -231 76 -197
<< metal1 >>
rect -88 231 -30 237
rect -88 197 -76 231
rect -42 197 -30 231
rect -88 191 -30 197
rect 30 231 88 237
rect 30 197 42 231
rect 76 197 88 231
rect 30 191 88 197
rect -141 138 -95 150
rect -141 -138 -135 138
rect -101 -138 -95 138
rect -141 -150 -95 -138
rect -23 138 23 150
rect -23 -138 -17 138
rect 17 -138 23 138
rect -23 -150 23 -138
rect 95 138 141 150
rect 95 -138 101 138
rect 135 -138 141 138
rect 95 -150 141 -138
rect -88 -197 -30 -191
rect -88 -231 -76 -197
rect -42 -231 -30 -197
rect -88 -237 -30 -231
rect 30 -197 88 -191
rect 30 -231 42 -197
rect 76 -231 88 -197
rect 30 -237 88 -231
<< properties >>
string FIXED_BBOX -232 -316 232 316
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.5 l 0.3 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

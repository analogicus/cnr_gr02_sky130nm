magic
tech sky130B
magscale 1 2
timestamp 1713519087
<< nwell >>
rect -226 -484 226 484
<< pmos >>
rect -30 -336 30 264
<< pdiff >>
rect -88 252 -30 264
rect -88 -324 -76 252
rect -42 -324 -30 252
rect -88 -336 -30 -324
rect 30 252 88 264
rect 30 -324 42 252
rect 76 -324 88 252
rect 30 -336 88 -324
<< pdiffc >>
rect -76 -324 -42 252
rect 42 -324 76 252
<< nsubdiff >>
rect -156 414 -94 448
rect 94 414 156 448
rect -156 -448 -94 -414
rect 94 -448 156 -414
<< nsubdiffcont >>
rect -94 414 94 448
rect -94 -448 94 -414
<< poly >>
rect -197 -375 -149 355
rect -33 345 33 361
rect -33 311 -17 345
rect 17 311 33 345
rect -33 295 33 311
rect -30 264 30 295
rect -30 -362 30 -336
rect 153 -373 201 357
<< polycont >>
rect -17 311 17 345
<< locali >>
rect -110 414 -94 448
rect 94 414 110 448
rect -33 311 -17 345
rect 17 311 33 345
rect -76 252 -42 268
rect -76 -340 -42 -324
rect 42 252 76 268
rect 42 -340 76 -324
rect -110 -448 -94 -414
rect 94 -448 110 -414
<< viali >>
rect -17 311 17 345
rect -76 -324 -42 252
rect 42 -324 76 252
<< metal1 >>
rect -39 345 39 359
rect -39 311 -17 345
rect 17 311 39 345
rect -39 299 39 311
rect -82 252 -36 264
rect -82 -324 -76 252
rect -42 -324 -36 252
rect -82 -336 -36 -324
rect 36 252 82 264
rect 36 -324 42 252
rect 76 -324 82 252
rect 36 -336 82 -324
<< properties >>
string FIXED_BBOX -173 -431 173 431
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3 l .3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/RPLY_EX0_lpe.spi
#else
.include ../../../work/xsch/RPLY_EX0.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6 keepopinfo noopiter gminsteps=5

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p


*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD  0  dc 1.8

*-----------------------------------------------------------------
* To test OTA
*-----------------------------------------------------------------
*Rin1	in1	vcm1	100
*Rin2	in2	vcm2	100

*vcm1	vcm1	0	dc	.7
*vcm2	vcm2	0	dc	.7
*vin	in1	in2	sin(0	10m	1K)

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VDD VSS RPLY_EX0

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.save v(VDD) v(VSS) v(in1) v(in2) v(xdut.VRO0) v(xdut.vbjt1) v(xdut.vo) v(xdut.VBJT2) v(xdut.vro)

#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

save @m.xdut.xm4.msky130_fd_pr__pfet_01v8[id]
+ @m.xdut.xm4.msky130_fd_pr__pfet_01v8[vgs]
+ @m.xdut.xm4.msky130_fd_pr__pfet_01v8[vds]
+ @m.xdut.xm4.msky130_fd_pr__pfet_01v8[vth]
+ @m.xdut.xm1.msky130_fd_pr__pfet_01v8[vgs]
+ @m.xdut.xm1.msky130_fd_pr__pfet_01v8[vth]
+ @m.xdut.xm1.msky130_fd_pr__pfet_01v8[vds]
+ @m.xdut.xm1.msky130_fd_pr__pfet_01v8[id]
+ @m.xdut.xm2.msky130_fd_pr__pfet_01v8[vgs]
+ @m.xdut.xm2.msky130_fd_pr__pfet_01v8[vth]
+ @m.xdut.xm2.msky130_fd_pr__pfet_01v8[vds]
+ @m.xdut.xm2.msky130_fd_pr__pfet_01v8[id]
+ @m.xdut.xm3.msky130_fd_pr__pfet_01v8[vgs]
+ @m.xdut.xm3.msky130_fd_pr__pfet_01v8[vth]
+ @m.xdut.xm3.msky130_fd_pr__pfet_01v8[vds]
+ @m.xdut.xm3.msky130_fd_pr__pfet_01v8[id]
+ @m.xdut.xm9.msky130_fd_pr__pfet_01v8[id]
+ @m.xdut.xm9.msky130_fd_pr__pfet_01v8[vgs]
+ @m.xdut.xm9.msky130_fd_pr__pfet_01v8[vds]
+ @m.xdut.xm9.msky130_fd_pr__pfet_01v8[vth]
+ @m.xdut.xm10.msky130_fd_pr__pfet_01v8[id]
+ @m.xdut.xm10.msky130_fd_pr__pfet_01v8[vgs]
+ @m.xdut.xm10.msky130_fd_pr__pfet_01v8[vds]
+ @m.xdut.xm10.msky130_fd_pr__pfet_01v8[vth]
+ @m.xdut.xm11.msky130_fd_pr__pfet_01v8[id]
+ @m.xdut.xm11.msky130_fd_pr__pfet_01v8[vgs]
+ @m.xdut.xm11.msky130_fd_pr__pfet_01v8[vds]
+ @m.xdut.xm11.msky130_fd_pr__pfet_01v8[vth]
+ @m.xdut.xm12.msky130_fd_pr__pfet_01v8[id]
+ @m.xdut.xm12.msky130_fd_pr__pfet_01v8[vgs]
+ @m.xdut.xm12.msky130_fd_pr__pfet_01v8[vds]
+ @m.xdut.xm12.msky130_fd_pr__pfet_01v8[vth]
+ @m.xdut.xm13.msky130_fd_pr__pfet_01v8[id]
+ @m.xdut.xm13.msky130_fd_pr__pfet_01v8[vgs]
+ @m.xdut.xm13.msky130_fd_pr__pfet_01v8[vds]
+ @m.xdut.xm13.msky130_fd_pr__pfet_01v8[vth]
+ @m.xdut.xm14.msky130_fd_pr__pfet_01v8[id]
+ @m.xdut.xm14.msky130_fd_pr__pfet_01v8[vgs]
+ @m.xdut.xm14.msky130_fd_pr__pfet_01v8[vds]
+ @m.xdut.xm14.msky130_fd_pr__pfet_01v8[vth]
+ @m.xdut.xm16.msky130_fd_pr__pfet_01v8[id]
+ @m.xdut.xm16.msky130_fd_pr__pfet_01v8[vgs]
+ @m.xdut.xm16.msky130_fd_pr__pfet_01v8[vds]
+ @m.xdut.xm16.msky130_fd_pr__pfet_01v8[vth]


+ @m.xdut.xm5.msky130_fd_pr__nfet_01v8[id]
+ @m.xdut.xm5.msky130_fd_pr__nfet_01v8[vgs]
+ @m.xdut.xm5.msky130_fd_pr__nfet_01v8[vds]
+ @m.xdut.xm5.msky130_fd_pr__nfet_01v8[vth]
+ @m.xdut.xm6.msky130_fd_pr__nfet_01v8[id]
+ @m.xdut.xm6.msky130_fd_pr__nfet_01v8[vgs]
+ @m.xdut.xm6.msky130_fd_pr__nfet_01v8[vds]
+ @m.xdut.xm6.msky130_fd_pr__nfet_01v8[vth]
+ @m.xdut.xm7.msky130_fd_pr__nfet_01v8[id]
+ @m.xdut.xm7.msky130_fd_pr__nfet_01v8[vgs]
+ @m.xdut.xm7.msky130_fd_pr__nfet_01v8[vds]
+ @m.xdut.xm8.msky130_fd_pr__nfet_01v8[id]
+ @m.xdut.xm8.msky130_fd_pr__nfet_01v8[vgs]
+ @m.xdut.xm8.msky130_fd_pr__nfet_01v8[vds]
+ @m.xdut.xm8.msky130_fd_pr__nfet_01v8[vth]



op


let vo=v(xdut.vo)
*let vbjt2=v(xdut.VBJT2)
let vref=v(xdut.vro)
let vbjt1=v(xdut.vbjt1)
let vro0=v(xdut.vro0)
let vdf=v(xdut.vbjt1)-v(xdut.vro0)


let i16 = @m.xdut.xm16.msky130_fd_pr__pfet_01v8[id]
let s16=@m.xdut.xm16.msky130_fd_pr__pfet_01v8[vds]-@m.xdut.xm16.msky130_fd_pr__pfet_01v8[vgs]+@m.xdut.xm16.msky130_fd_pr__pfet_01v8[vth]
let vgs16 = @m.xdut.xm16.msky130_fd_pr__pfet_01v8[vgs]
let vds16 = @m.xdut.xm16.msky130_fd_pr__pfet_01v8[vds]
let i4 = @m.xdut.xm4.msky130_fd_pr__pfet_01v8[id]
let s4=@m.xdut.xm4.msky130_fd_pr__pfet_01v8[vds]-@m.xdut.xm4.msky130_fd_pr__pfet_01v8[vgs]+@m.xdut.xm4.msky130_fd_pr__pfet_01v8[vth]
let vgs4 = @m.xdut.xm4.msky130_fd_pr__pfet_01v8[vgs]
let vds4 = @m.xdut.xm4.msky130_fd_pr__pfet_01v8[vds]
let i3 = @m.xdut.xm3.msky130_fd_pr__pfet_01v8[id]
let s3=@m.xdut.xm3.msky130_fd_pr__pfet_01v8[vds]-@m.xdut.xm3.msky130_fd_pr__pfet_01v8[vgs]+@m.xdut.xm3.msky130_fd_pr__pfet_01v8[vth]
let vgs3 = @m.xdut.xm3.msky130_fd_pr__pfet_01v8[vgs]
let vds3 = @m.xdut.xm3.msky130_fd_pr__pfet_01v8[vds]
let i1 = @m.xdut.xm1.msky130_fd_pr__pfet_01v8[id]
let vgs1 = @m.xdut.xm1.msky130_fd_pr__pfet_01v8[vgs]
let vds1 = @m.xdut.xm1.msky130_fd_pr__pfet_01v8[vds]
let s1=@m.xdut.xm1.msky130_fd_pr__pfet_01v8[vds]-@m.xdut.xm1.msky130_fd_pr__pfet_01v8[vgs]+@m.xdut.xm1.msky130_fd_pr__pfet_01v8[vth]
let i2 = @m.xdut.xm2.msky130_fd_pr__pfet_01v8[id]
let vgs2 = @m.xdut.xm2.msky130_fd_pr__pfet_01v8[vgs]
let vds2 = @m.xdut.xm2.msky130_fd_pr__pfet_01v8[vds]
let s2=@m.xdut.xm2.msky130_fd_pr__pfet_01v8[vds]-@m.xdut.xm2.msky130_fd_pr__pfet_01v8[vgs]+@m.xdut.xm2.msky130_fd_pr__pfet_01v8[vth]
let s9=@m.xdut.xm9.msky130_fd_pr__pfet_01v8[vds]-@m.xdut.xm9.msky130_fd_pr__pfet_01v8[vgs]+@m.xdut.xm9.msky130_fd_pr__pfet_01v8[vth]
let i9=@m.xdut.xm9.msky130_fd_pr__pfet_01v8[id]
let vgs9=@m.xdut.xm9.msky130_fd_pr__pfet_01v8[vgs]
let vds9=@m.xdut.xm9.msky130_fd_pr__pfet_01v8[vds]
let s10=@m.xdut.xm10.msky130_fd_pr__pfet_01v8[vds]-@m.xdut.xm10.msky130_fd_pr__pfet_01v8[vgs]+@m.xdut.xm10.msky130_fd_pr__pfet_01v8[vth]
let vgs10=@m.xdut.xm10.msky130_fd_pr__pfet_01v8[vgs]
let vds10=@m.xdut.xm10.msky130_fd_pr__pfet_01v8[vds]
let i10 = @m.xdut.xm10.msky130_fd_pr__pfet_01v8[id]
let i11 = @m.xdut.xm11.msky130_fd_pr__pfet_01v8[id]
let s11= @m.xdut.xm11.msky130_fd_pr__pfet_01v8[vds]-@m.xdut.xm11.msky130_fd_pr__pfet_01v8[vgs]+@m.xdut.xm11.msky130_fd_pr__pfet_01v8[vth]
let vgs11 = @m.xdut.xm11.msky130_fd_pr__pfet_01v8[vgs]
let vds11 = @m.xdut.xm11.msky130_fd_pr__pfet_01v8[vds]
let i12 = @m.xdut.xm12.msky130_fd_pr__pfet_01v8[id]
let s12 = @m.xdut.xm12.msky130_fd_pr__pfet_01v8[vds]-@m.xdut.xm12.msky130_fd_pr__pfet_01v8[vgs]+@m.xdut.xm12.msky130_fd_pr__pfet_01v8[vth]
let vgs12 = @m.xdut.xm12.msky130_fd_pr__pfet_01v8[vgs]
let vds12 = @m.xdut.xm12.msky130_fd_pr__pfet_01v8[vds]
let i13 = @m.xdut.xm13.msky130_fd_pr__pfet_01v8[id]
let s13 = @m.xdut.xm13.msky130_fd_pr__pfet_01v8[vds]-@m.xdut.xm13.msky130_fd_pr__pfet_01v8[vgs]+@m.xdut.xm13.msky130_fd_pr__pfet_01v8[vth]
let vgs13 = @m.xdut.xm13.msky130_fd_pr__pfet_01v8[vgs]
let vds13 = @m.xdut.xm13.msky130_fd_pr__pfet_01v8[vds]
let i14 = @m.xdut.xm14.msky130_fd_pr__pfet_01v8[id]
let vgs14 = @m.xdut.xm14.msky130_fd_pr__pfet_01v8[vgs]
let vds14 = @m.xdut.xm14.msky130_fd_pr__pfet_01v8[vds]
let s14 = @m.xdut.xm14.msky130_fd_pr__pfet_01v8[vds]-@m.xdut.xm14.msky130_fd_pr__pfet_01v8[vgs]+@m.xdut.xm14.msky130_fd_pr__pfet_01v8[vth]



let i7 = @m.xdut.xm7.msky130_fd_pr__nfet_01v8[id]
let s7=@m.xdut.xm7.msky130_fd_pr__nfet_01v8[vds]-@m.xdut.xm7.msky130_fd_pr__nfet_01v8[vgs]+@m.xdut.xm7.msky130_fd_pr__nfet_01v8[vth]
let vgs7 = @m.xdut.xm7.msky130_fd_pr__nfet_01v8[vgs]
let vds7 = @m.xdut.xm7.msky130_fd_pr__nfet_01v8[vds]
let i8 = @m.xdut.xm8.msky130_fd_pr__nfet_01v8[id]
let s8=@m.xdut.xm8.msky130_fd_pr__nfet_01v8[vds]-@m.xdut.xm8.msky130_fd_pr__nfet_01v8[vgs]+@m.xdut.xm8.msky130_fd_pr__nfet_01v8[vth]
let vgs8 = @m.xdut.xm8.msky130_fd_pr__nfet_01v8[vgs]
let vds8 = @m.xdut.xm8.msky130_fd_pr__nfet_01v8[vds]
let i5 = @m.xdut.xm5.msky130_fd_pr__nfet_01v8[id]
let s5 = @m.xdut.xm5.msky130_fd_pr__nfet_01v8[vds]-@m.xdut.xm5.msky130_fd_pr__nfet_01v8[vgs]+@m.xdut.xm5.msky130_fd_pr__nfet_01v8[vth]
let vgs5 = @m.xdut.xm5.msky130_fd_pr__nfet_01v8[vgs]
let vds5 = @m.xdut.xm5.msky130_fd_pr__nfet_01v8[vds]
let i6 = @m.xdut.xm6.msky130_fd_pr__nfet_01v8[id]
let s6 = @m.xdut.xm6.msky130_fd_pr__nfet_01v8[vds]-@m.xdut.xm6.msky130_fd_pr__nfet_01v8[vgs]+@m.xdut.xm6.msky130_fd_pr__nfet_01v8[vth]
let vgs6 = @m.xdut.xm6.msky130_fd_pr__nfet_01v8[vgs]
let vds6 = @m.xdut.xm6.msky130_fd_pr__nfet_01v8[vds]



write
quit
#endif

.endc

.end

*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_GR02_lpe.spi
#else
.include ../../../work/xsch/CNR_GR02.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TEMP=40 GMIN=1e-15 reltol=1e-6 abstol=1e-6 keepopinfo noopiter gminsteps=5

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS VSS 0 dc 0
VDD_1V8 VDD_1V8 0 dc 1.8
Vrst rst 0 pwl 0 1.8 10u 1.8 10.01u 0
Vopamp LPO LPI dc 0
*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VDD_1V8 VSS rst VO LPO LPI CNR_GR02

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

.save all

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
set file = "tdiff.txt"
unset askquit

optran 0 0 0 100n 20u 0
* -40 -30 -20 -10 0 10 20 30 40 50 60 70 80 90 100 110 120
foreach vtemp 27
  option temp=$vtemp
  tran 100n 175u
  meas tran tdiff_$vtemp TRIG V(rst) VAL=0.5 FALL=1 TARG V(xdut.vop) VAL=.5 FALL=1 >> $file
  write {cicname}_$vtemp
end

* Checks
*let vd2branch = v(xdut.D2_Branch)
*let vref=v(xdut.D2_branch)-v(xdut.D2)
*let vd= v(xdut.D1)-v(xdut.D2_Branch) 
*let lpo=v(LPO)

write
quit
#endif

.endc

.end

magic
tech sky130B
magscale 1 2
timestamp 1713258222
<< pwell >>
rect -201 -1224 201 1224
<< psubdiff >>
rect -165 1154 -69 1188
rect 69 1154 165 1188
rect -165 1092 -131 1154
rect 131 1092 165 1154
rect -165 -1154 -131 -1092
rect 131 -1154 165 -1092
rect -165 -1188 -69 -1154
rect 69 -1188 165 -1154
<< psubdiffcont >>
rect -69 1154 69 1188
rect -165 -1092 -131 1092
rect 131 -1092 165 1092
rect -69 -1188 69 -1154
<< xpolycontact >>
rect -35 626 35 1058
rect -35 -1058 35 -626
<< ppolyres >>
rect -35 -626 35 626
<< locali >>
rect -165 1154 -69 1188
rect 69 1154 165 1188
rect -165 1092 -131 1154
rect 131 1092 165 1154
rect -165 -1154 -131 -1092
rect 131 -1154 165 -1092
rect -165 -1188 -69 -1154
rect 69 -1188 165 -1154
<< viali >>
rect -19 643 19 1040
rect -19 -1040 19 -643
<< metal1 >>
rect -25 1040 25 1052
rect -25 643 -19 1040
rect 19 643 25 1040
rect -25 631 25 643
rect -25 -643 25 -631
rect -25 -1040 -19 -643
rect 19 -1040 25 -643
rect -25 -1052 25 -1040
<< properties >>
string FIXED_BBOX -148 -1171 148 1171
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.35 l 6.42 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 6.979k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

magic
tech sky130B
magscale 1 2
timestamp 1713258222
<< nwell >>
rect -1825 -969 1825 969
<< pmos >>
rect -1629 -750 -29 750
rect 29 -750 1629 750
<< pdiff >>
rect -1687 738 -1629 750
rect -1687 -738 -1675 738
rect -1641 -738 -1629 738
rect -1687 -750 -1629 -738
rect -29 738 29 750
rect -29 -738 -17 738
rect 17 -738 29 738
rect -29 -750 29 -738
rect 1629 738 1687 750
rect 1629 -738 1641 738
rect 1675 -738 1687 738
rect 1629 -750 1687 -738
<< pdiffc >>
rect -1675 -738 -1641 738
rect -17 -738 17 738
rect 1641 -738 1675 738
<< nsubdiff >>
rect -1789 899 -1693 933
rect 1693 899 1789 933
rect -1789 837 -1755 899
rect 1755 837 1789 899
rect -1789 -899 -1755 -837
rect 1755 -899 1789 -837
rect -1789 -933 -1693 -899
rect 1693 -933 1789 -899
<< nsubdiffcont >>
rect -1693 899 1693 933
rect -1789 -837 -1755 837
rect 1755 -837 1789 837
rect -1693 -933 1693 -899
<< poly >>
rect -1629 831 -29 847
rect -1629 797 -1613 831
rect -45 797 -29 831
rect -1629 750 -29 797
rect 29 831 1629 847
rect 29 797 45 831
rect 1613 797 1629 831
rect 29 750 1629 797
rect -1629 -797 -29 -750
rect -1629 -831 -1613 -797
rect -45 -831 -29 -797
rect -1629 -847 -29 -831
rect 29 -797 1629 -750
rect 29 -831 45 -797
rect 1613 -831 1629 -797
rect 29 -847 1629 -831
<< polycont >>
rect -1613 797 -45 831
rect 45 797 1613 831
rect -1613 -831 -45 -797
rect 45 -831 1613 -797
<< locali >>
rect -1789 899 -1693 933
rect 1693 899 1789 933
rect -1789 837 -1755 899
rect 1755 837 1789 899
rect -1629 797 -1613 831
rect -45 797 -29 831
rect 29 797 45 831
rect 1613 797 1629 831
rect -1675 738 -1641 754
rect -1675 -754 -1641 -738
rect -17 738 17 754
rect -17 -754 17 -738
rect 1641 738 1675 754
rect 1641 -754 1675 -738
rect -1629 -831 -1613 -797
rect -45 -831 -29 -797
rect 29 -831 45 -797
rect 1613 -831 1629 -797
rect -1789 -899 -1755 -837
rect 1755 -899 1789 -837
rect -1789 -933 -1693 -899
rect 1693 -933 1789 -899
<< viali >>
rect -1613 797 -45 831
rect 45 797 1613 831
rect -1675 -738 -1641 738
rect -17 -738 17 738
rect 1641 -738 1675 738
rect -1613 -831 -45 -797
rect 45 -831 1613 -797
<< metal1 >>
rect -1625 831 -33 837
rect -1625 797 -1613 831
rect -45 797 -33 831
rect -1625 791 -33 797
rect 33 831 1625 837
rect 33 797 45 831
rect 1613 797 1625 831
rect 33 791 1625 797
rect -1681 738 -1635 750
rect -1681 -738 -1675 738
rect -1641 -738 -1635 738
rect -1681 -750 -1635 -738
rect -23 738 23 750
rect -23 -738 -17 738
rect 17 -738 23 738
rect -23 -750 23 -738
rect 1635 738 1681 750
rect 1635 -738 1641 738
rect 1675 -738 1681 738
rect 1635 -750 1681 -738
rect -1625 -797 -33 -791
rect -1625 -831 -1613 -797
rect -45 -831 -33 -797
rect -1625 -837 -33 -831
rect 33 -797 1625 -791
rect 33 -831 45 -797
rect 1613 -831 1625 -797
rect 33 -837 1625 -831
<< properties >>
string FIXED_BBOX -1772 -916 1772 916
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 7.5 l 8.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

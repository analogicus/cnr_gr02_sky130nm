** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/OTA_SKY130NM/TB_OTA.sch
**.subckt TB_OTA
V2 VIP GND 0.9
C1 VIN GND 1p m=1
V1 net1 GND 1.8
x1 net1 net2 net2 VIN VIN VIP GND OTA
**** begin user architecture code



* ngspice commands
.include corner.spi



**** end user architecture code
**.ends

* expanding   symbol:  OTA_SKY130NM/OTA.sym # of pins=7
** sym_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/OTA_SKY130NM/OTA.sym
** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/OTA_SKY130NM/OTA.sch
.subckt OTA VDD_1V8 LPO LPI VO VIN VIP VSS
*.ipin VSS
*.ipin VDD_1V8
*.ipin VIN
*.ipin VIP
*.opin VO
*.opin LPO
*.ipin LPI
R2 LPI VO sky130_fd_pr__res_generic_m1 W=1 L=1 m=1
x2 p5 VIN p1 p1 CNRATR_NCH_8C2F0
x3 p6 VIP p1 p1 CNRATR_NCH_8C2F0
x7 p6 p6 VDD_1V8 VDD_1V8 CNRATR_PCH_8C2F0
x9 LPO p6 VDD_1V8 VDD_1V8 CNRATR_PCH_12C4F0
x8 p3 p5 VDD_1V8 VDD_1V8 CNRATR_PCH_8C4F0
x5 p5 p5 VDD_1V8 VDD_1V8 CNRATR_PCH_8C2F0
x6 p1 p2 VSS VSS CNRATR_NCH_8C2F0
x1 p2 p2 VSS VSS CNRATR_NCH_8C2F0
x10 p3 p3 VSS VSS CNRATR_NCH_4C8F0
x11 LPO p3 VSS VSS CNRATR_NCH_12C12F0
I0 VDD_1V8 p2 3u
.ends


* expanding   symbol:  ../CNR_ATR_SKY130NM/CNRATR_NCH_8C2F0.sym # of pins=4
** sym_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_8C2F0.sym
** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_8C2F0.sch
.subckt CNRATR_NCH_8C2F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.54 W=7.68 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  ../CNR_ATR_SKY130NM/CNRATR_PCH_8C2F0.sym # of pins=4
** sym_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_8C2F0.sym
** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_8C2F0.sch
.subckt CNRATR_PCH_8C2F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.54 W=7.68 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  ../CNR_ATR_SKY130NM/CNRATR_PCH_12C4F0.sym # of pins=4
** sym_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_12C4F0.sym
** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_12C4F0.sch
.subckt CNRATR_PCH_12C4F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=1.26 W=11.52 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  ../CNR_ATR_SKY130NM/CNRATR_PCH_8C4F0.sym # of pins=4
** sym_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_8C4F0.sym
** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_8C4F0.sch
.subckt CNRATR_PCH_8C4F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=1.26 W=7.68 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  ../CNR_ATR_SKY130NM/CNRATR_NCH_4C8F0.sym # of pins=4
** sym_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_4C8F0.sym
** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_4C8F0.sch
.subckt CNRATR_NCH_4C8F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=2.7 W=3.84 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  ../CNR_ATR_SKY130NM/CNRATR_NCH_12C12F0.sym # of pins=4
** sym_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_12C12F0.sym
** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_12C12F0.sch
.subckt CNRATR_NCH_12C12F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=4.14 W=11.52 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end

magic
tech sky130B
timestamp 1713476340
<< pwell >>
rect -100 -873 100 873
<< psubdiff >>
rect -82 807 -65 838
rect -82 -838 -65 -807
<< psubdiffcont >>
rect -82 -807 -65 807
<< xpolycontact >>
rect -17 574 17 790
rect -17 -790 17 -574
<< ppolyres >>
rect -17 -574 17 574
<< locali >>
rect -82 807 -65 838
rect -82 -838 -65 -807
<< viali >>
rect -9 583 9 781
rect -9 -781 9 -583
<< metal1 >>
rect -12 781 12 787
rect -12 583 -9 781
rect 9 583 12 781
rect -12 577 12 583
rect -12 -583 12 -577
rect -12 -781 -9 -583
rect 9 -781 12 -583
rect -12 -787 12 -781
<< properties >>
string FIXED_BBOX -74 -847 74 847
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.35 l 11.65 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 11.758k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

magic
tech sky130B
magscale 1 2
timestamp 1713313793
<< locali >>
rect -6110 910 -4580 1050
rect -6110 830 -5920 910
rect -4770 830 -4580 910
rect -4540 870 -4250 1050
rect -4210 910 -2680 1050
rect -5960 440 -5680 670
rect -6000 -190 -5680 40
rect -5024 28 -4960 410
rect -5267 -109 -4965 -39
rect -4425 -44 -4354 870
rect -4210 830 -4020 910
rect -2870 830 -2680 910
rect -4120 410 -3800 640
rect -3365 493 -2927 559
rect -4426 -104 -4420 -44
rect -4360 -104 -4354 -44
rect -4426 -110 -4354 -104
rect -4120 -190 -3800 40
rect -3540 -106 -3536 -42
rect -3464 -106 -3058 -42
rect -6010 -800 -5690 -570
rect -5450 -710 -5446 -640
rect -5374 -710 -5370 -640
rect -5155 -705 -4966 -636
rect -6030 -1400 -5684 -1170
rect -5155 -1240 -5086 -705
rect -4100 -800 -3780 -570
rect -3124 -712 -3059 -203
rect -5309 -1309 -5086 -1240
rect -4100 -1400 -3780 -1170
rect -2993 -1247 -2927 493
rect -3123 -1313 -2927 -1247
rect -4525 -1691 -3175 -1685
rect -4525 -1749 -4519 -1691
rect -4461 -1749 -3175 -1691
rect -4525 -1755 -3175 -1749
rect -6030 -1990 -5684 -1760
rect -4392 -1834 -4328 -1828
rect -5285 -1910 -4965 -1839
rect -4392 -1886 -4386 -1834
rect -4334 -1886 -4328 -1834
rect -6030 -2590 -5684 -2360
rect -5023 -2431 -4961 -2005
rect -5440 -2510 -5109 -2446
rect -4392 -2448 -4328 -1886
rect -4130 -2280 -3794 -2050
rect -3245 -2135 -3175 -1755
rect -3555 -2205 -3175 -2135
rect -3118 -2443 -3065 -2309
rect -5172 -2786 -5109 -2510
rect -4392 -2512 -4088 -2448
rect -3193 -2496 -3065 -2443
rect -5861 -2848 -5108 -2786
rect -4392 -2848 -4329 -2672
rect -5861 -2849 -4329 -2848
rect -5861 -2980 -5798 -2849
rect -5172 -2911 -4329 -2849
rect -4140 -2880 -3774 -2650
rect -6110 -3110 -5600 -2980
rect -5460 -3039 -4950 -2980
rect -5460 -3080 -5247 -3039
rect -5206 -3080 -4950 -3039
rect -5460 -3110 -4950 -3080
rect -4840 -3034 -4330 -2980
rect -4840 -3083 -4684 -3034
rect -4635 -3083 -4330 -3034
rect -4840 -3110 -4330 -3083
rect -3122 -3029 -3061 -2905
<< viali >>
rect -5441 489 -5374 556
rect -5440 -110 -5380 -50
rect -3540 493 -3481 552
rect -4420 -104 -4360 -44
rect -3536 -110 -3464 -38
rect -5446 -710 -5374 -638
rect -5440 -1302 -5376 -1238
rect -3540 -710 -3476 -646
rect -5010 -1330 -4970 -1250
rect -3535 -1296 -3484 -1245
rect -4519 -1749 -4461 -1691
rect -5434 -1906 -5382 -1854
rect -4386 -1886 -4334 -1834
rect -5013 -2484 -4966 -2437
rect -3246 -2496 -3193 -2443
rect -4392 -2672 -4329 -2609
rect -3540 -2810 -3481 -2738
rect -5247 -3080 -5206 -3039
rect -4684 -3083 -4635 -3034
rect -3122 -3090 -3061 -3029
<< metal1 >>
rect -5447 558 -5368 568
rect -5447 556 -3469 558
rect -5447 489 -5441 556
rect -5374 552 -3469 556
rect -5374 493 -3540 552
rect -3481 493 -3469 552
rect -5374 489 -3469 493
rect -5447 487 -3469 489
rect -5447 477 -5368 487
rect -4426 -38 -4354 -32
rect -3542 -38 -3458 -26
rect -5446 -50 -5374 -38
rect -5446 -110 -5440 -50
rect -5380 -110 -5374 -50
rect -5446 -340 -5374 -110
rect -4426 -44 -3536 -38
rect -4426 -104 -4420 -44
rect -4360 -104 -3536 -44
rect -4426 -110 -3536 -104
rect -3464 -110 -3458 -38
rect -4426 -116 -4354 -110
rect -3542 -122 -3458 -110
rect -5450 -410 -4820 -340
rect -5446 -632 -5374 -410
rect -5458 -638 -5362 -632
rect -5458 -710 -5446 -638
rect -5374 -710 -5362 -638
rect -5458 -716 -5362 -710
rect -5452 -1238 -5364 -1232
rect -5452 -1302 -5440 -1238
rect -5376 -1302 -5364 -1238
rect -5452 -1308 -5364 -1302
rect -5030 -1250 -4950 -1230
rect -4890 -1250 -4820 -410
rect -3546 -646 -3470 -634
rect -5440 -1854 -5376 -1308
rect -5030 -1330 -5010 -1250
rect -4970 -1320 -4820 -1250
rect -4970 -1330 -4950 -1320
rect -5030 -1340 -4950 -1330
rect -4890 -1685 -4820 -1320
rect -4392 -710 -3540 -646
rect -3476 -710 -3470 -646
rect -4890 -1691 -4449 -1685
rect -4890 -1749 -4519 -1691
rect -4461 -1749 -4449 -1691
rect -4890 -1755 -4449 -1749
rect -5440 -1906 -5434 -1854
rect -5382 -1906 -5376 -1854
rect -4392 -1834 -4328 -710
rect -3546 -722 -3470 -710
rect -3547 -1245 -3179 -1239
rect -3547 -1296 -3535 -1245
rect -3484 -1296 -3179 -1245
rect -3547 -1302 -3179 -1296
rect -4392 -1886 -4386 -1834
rect -4334 -1886 -4328 -1834
rect -4392 -1898 -4328 -1886
rect -5440 -1918 -5376 -1906
rect -3242 -1959 -3179 -1302
rect -4391 -2022 -3179 -1959
rect -5019 -2437 -4960 -2425
rect -5019 -2484 -5013 -2437
rect -4966 -2484 -4960 -2437
rect -5019 -2744 -4960 -2484
rect -4391 -2603 -4328 -2022
rect -3258 -2443 -3181 -2437
rect -3258 -2496 -3246 -2443
rect -3193 -2496 -3181 -2443
rect -3258 -2502 -3181 -2496
rect -4404 -2609 -4317 -2603
rect -4404 -2672 -4392 -2609
rect -4329 -2672 -4317 -2609
rect -4404 -2678 -4317 -2672
rect -3546 -2738 -3475 -2726
rect -3546 -2744 -3540 -2738
rect -5019 -2803 -3540 -2744
rect -3546 -2810 -3540 -2803
rect -3481 -2810 -3475 -2738
rect -3546 -2822 -3475 -2810
rect -3245 -2863 -3192 -2502
rect -5253 -2916 -3192 -2863
rect -5253 -3039 -5200 -2916
rect -3134 -3028 -3049 -3023
rect -5253 -3080 -5247 -3039
rect -5206 -3080 -5200 -3039
rect -5253 -3092 -5200 -3080
rect -4696 -3029 -3049 -3028
rect -4696 -3034 -3122 -3029
rect -4696 -3083 -4684 -3034
rect -4635 -3083 -3122 -3034
rect -4696 -3089 -3122 -3083
rect -3134 -3090 -3122 -3089
rect -3061 -3090 -3049 -3029
rect -3134 -3096 -3049 -3090
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713296683
transform 1 0 -4116 0 1 224
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_1
timestamp 1713296683
transform 1 0 -4116 0 1 -376
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_2
timestamp 1713296683
transform 1 0 -4116 0 1 -3076
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_3
timestamp 1713296683
transform 1 0 -4116 0 1 -976
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_4
timestamp 1713296683
transform 1 0 -4116 0 1 -2476
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_5
timestamp 1713296683
transform 1 0 -4116 0 1 -1576
box -184 -124 1528 728
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 -6016 0 1 224
box -184 -124 1528 728
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_1
timestamp 1695852000
transform 1 0 -6016 0 1 -376
box -184 -124 1528 728
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_2
timestamp 1695852000
transform 1 0 -6016 0 1 -976
box -184 -124 1528 728
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_3
timestamp 1695852000
transform 1 0 -6016 0 1 -1576
box -184 -124 1528 728
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_4
timestamp 1695852000
transform 1 0 -6016 0 1 -2176
box -184 -124 1528 728
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_5
timestamp 1695852000
transform 1 0 -6016 0 1 -2776
box -184 -124 1528 728
<< labels >>
flabel locali -5670 930 -5000 1030 0 FreeSans 400 0 0 0 VDD
port 1 nsew
flabel locali -3850 920 -3030 1030 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel locali -4520 880 -4270 1040 0 FreeSans 400 0 0 0 I_BIAS
port 4 nsew
flabel locali -5420 -3100 -4990 -2990 0 FreeSans 400 0 0 0 VIN
port 5 nsew
flabel locali -4800 -3100 -4370 -2990 0 FreeSans 400 0 0 0 VIP
port 6 nsew
flabel locali -6070 -3100 -5640 -2990 0 FreeSans 400 0 0 0 VO
port 7 nsew
<< end >>

magic
tech sky130B
magscale 1 2
timestamp 1713518785
<< pwell >>
rect -496 -379 496 379
<< nmos >>
rect -300 -231 300 169
<< ndiff >>
rect -358 157 -300 169
rect -358 -219 -346 157
rect -312 -219 -300 157
rect -358 -231 -300 -219
rect 300 157 358 169
rect 300 -219 312 157
rect 346 -219 358 157
rect 300 -231 358 -219
<< ndiffc >>
rect -346 -219 -312 157
rect 312 -219 346 157
<< psubdiff >>
rect -426 309 -364 343
rect 364 309 426 343
rect -426 -343 -364 -309
rect 364 -343 426 -309
<< psubdiffcont >>
rect -364 309 364 343
rect -364 -343 364 -309
<< poly >>
rect -473 -264 -417 246
rect -300 241 300 257
rect -300 207 -284 241
rect 284 207 300 241
rect -300 169 300 207
rect -300 -257 300 -231
rect 415 -248 471 262
<< polycont >>
rect -284 207 284 241
<< locali >>
rect -380 309 -364 343
rect 364 309 380 343
rect -300 207 -284 241
rect 284 207 300 241
rect -346 157 -312 173
rect -346 -235 -312 -219
rect 312 157 346 173
rect 312 -235 346 -219
rect -380 -343 -364 -309
rect 364 -343 380 -309
<< viali >>
rect -284 207 284 241
rect -346 -219 -312 157
rect 312 -219 346 157
<< metal1 >>
rect -296 241 296 247
rect -296 207 -284 241
rect 284 207 296 241
rect -296 201 296 207
rect -352 157 -306 169
rect -352 -219 -346 157
rect -312 -219 -306 157
rect -352 -231 -306 -219
rect 306 157 352 169
rect 306 -219 312 157
rect 346 -219 352 157
rect 306 -231 352 -219
<< properties >>
string FIXED_BBOX -443 -326 443 326
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

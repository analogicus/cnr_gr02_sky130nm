magic
tech sky130B
magscale 1 2
timestamp 1713555407
<< pwell >>
rect -201 -1237 201 1237
<< psubdiff >>
rect -165 1167 -69 1201
rect 69 1167 165 1201
rect -165 1105 -131 1167
rect 131 1105 165 1167
rect -165 -1167 -131 -1105
rect 131 -1167 165 -1105
rect -165 -1201 -69 -1167
rect 69 -1201 165 -1167
<< psubdiffcont >>
rect -69 1167 69 1201
rect -165 -1105 -131 1105
rect 131 -1105 165 1105
rect -69 -1201 69 -1167
<< xpolycontact >>
rect -35 639 35 1071
rect -35 -1071 35 -639
<< ppolyres >>
rect -35 -639 35 639
<< locali >>
rect -165 1167 -69 1201
rect 69 1167 165 1201
rect -165 1105 -131 1167
rect 131 1105 165 1167
rect -165 -1167 -131 -1105
rect 131 -1167 165 -1105
rect -165 -1201 -69 -1167
rect 69 -1201 165 -1167
<< viali >>
rect -19 656 19 1053
rect -19 -1053 19 -656
<< metal1 >>
rect -25 1053 25 1065
rect -25 656 -19 1053
rect 19 656 25 1053
rect -25 644 25 656
rect -25 -656 25 -644
rect -25 -1053 -19 -656
rect 19 -1053 25 -656
rect -25 -1065 25 -1053
<< properties >>
string FIXED_BBOX -148 -1184 148 1184
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 6.55 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 7.098k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

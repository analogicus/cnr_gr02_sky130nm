** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/OTA_SKY130NM/OTA.sch
.subckt OTA VSS VDD_1V8 LPI VIP LPO
*.ipin VSS
*.ipin VDD_1V8
*.ipin LPI
*.ipin VIP
*.opin LPO
x2 net3 LPI net1 net1 CNRATR_NCH_4C2F0
x3 net2 VIP net1 net1 CNRATR_NCH_4C2F0
x7 net2 net2 VDD_1V8 VDD_1V8 CNRATR_PCH_4C2F0
x9 net4 net2 VDD_1V8 VDD_1V8 CNRATR_PCH_4C2F0
x8 net5 net3 VDD_1V8 VDD_1V8 CNRATR_PCH_4C2F0
x5 net3 net3 VDD_1V8 VDD_1V8 CNRATR_PCH_4C2F0
x6 net1 net6 VSS VSS CNRATR_NCH_4C2F0
x1 net6 net6 VSS VSS CNRATR_NCH_4C2F0
x10 net5 net5 VSS VSS CNRATR_NCH_4C2F0
x11 net4 net5 VSS VSS CNRATR_NCH_4C2F0
I0 VDD_1V8 net6 5u
x12 net3 net2 VDD_1V8 VDD_1V8 CNRATR_PCH_2C2F0
x13 net2 net3 VDD_1V8 VDD_1V8 CNRATR_PCH_2C2F0
C1 LPO VSS 1p m=1
R1 net4 LPO 100k m=1
.ends

* expanding   symbol:  ../CNR_ATR_SKY130NM/CNRATR_NCH_4C2F0.sym # of pins=4
** sym_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_4C2F0.sym
** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_4C2F0.sch
.subckt CNRATR_NCH_4C2F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.54 W=3.84 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  ../CNR_ATR_SKY130NM/CNRATR_PCH_4C2F0.sym # of pins=4
** sym_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_4C2F0.sym
** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_4C2F0.sch
.subckt CNRATR_PCH_4C2F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.54 W=3.84 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  ../CNR_ATR_SKY130NM/CNRATR_PCH_2C2F0.sym # of pins=4
** sym_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_2C2F0.sym
** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_2C2F0.sch
.subckt CNRATR_PCH_2C2F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.54 W=1.92 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end

magic
tech sky130B
magscale 1 2
timestamp 1713258222
<< nwell >>
rect -425 -269 425 269
<< pmos >>
rect -229 -50 -29 50
rect 29 -50 229 50
<< pdiff >>
rect -287 38 -229 50
rect -287 -38 -275 38
rect -241 -38 -229 38
rect -287 -50 -229 -38
rect -29 38 29 50
rect -29 -38 -17 38
rect 17 -38 29 38
rect -29 -50 29 -38
rect 229 38 287 50
rect 229 -38 241 38
rect 275 -38 287 38
rect 229 -50 287 -38
<< pdiffc >>
rect -275 -38 -241 38
rect -17 -38 17 38
rect 241 -38 275 38
<< nsubdiff >>
rect -389 199 -293 233
rect 293 199 389 233
rect -389 137 -355 199
rect 355 137 389 199
rect -389 -199 -355 -137
rect 355 -199 389 -137
rect -389 -233 -293 -199
rect 293 -233 389 -199
<< nsubdiffcont >>
rect -293 199 293 233
rect -389 -137 -355 137
rect 355 -137 389 137
rect -293 -233 293 -199
<< poly >>
rect -229 131 -29 147
rect -229 97 -213 131
rect -45 97 -29 131
rect -229 50 -29 97
rect 29 131 229 147
rect 29 97 45 131
rect 213 97 229 131
rect 29 50 229 97
rect -229 -97 -29 -50
rect -229 -131 -213 -97
rect -45 -131 -29 -97
rect -229 -147 -29 -131
rect 29 -97 229 -50
rect 29 -131 45 -97
rect 213 -131 229 -97
rect 29 -147 229 -131
<< polycont >>
rect -213 97 -45 131
rect 45 97 213 131
rect -213 -131 -45 -97
rect 45 -131 213 -97
<< locali >>
rect -389 199 -293 233
rect 293 199 389 233
rect -389 137 -355 199
rect 355 137 389 199
rect -229 97 -213 131
rect -45 97 -29 131
rect 29 97 45 131
rect 213 97 229 131
rect -275 38 -241 54
rect -275 -54 -241 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 241 38 275 54
rect 241 -54 275 -38
rect -229 -131 -213 -97
rect -45 -131 -29 -97
rect 29 -131 45 -97
rect 213 -131 229 -97
rect -389 -199 -355 -137
rect 355 -199 389 -137
rect -389 -233 -293 -199
rect 293 -233 389 -199
<< viali >>
rect -213 97 -45 131
rect 45 97 213 131
rect -275 -38 -241 38
rect -17 -38 17 38
rect 241 -38 275 38
rect -213 -131 -45 -97
rect 45 -131 213 -97
<< metal1 >>
rect -225 131 -33 137
rect -225 97 -213 131
rect -45 97 -33 131
rect -225 91 -33 97
rect 33 131 225 137
rect 33 97 45 131
rect 213 97 225 131
rect 33 91 225 97
rect -281 38 -235 50
rect -281 -38 -275 38
rect -241 -38 -235 38
rect -281 -50 -235 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 235 38 281 50
rect 235 -38 241 38
rect 275 -38 281 38
rect 235 -50 281 -38
rect -225 -97 -33 -91
rect -225 -131 -213 -97
rect -45 -131 -33 -97
rect -225 -137 -33 -131
rect 33 -97 225 -91
rect 33 -131 45 -97
rect 213 -131 225 -97
rect 33 -137 225 -131
<< properties >>
string FIXED_BBOX -372 -216 372 216
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.5 l 1.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

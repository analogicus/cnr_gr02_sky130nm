magic
tech sky130B
magscale 1 2
timestamp 1713550659
<< nwell >>
rect 3960 3042 6445 4120
rect 9900 3166 12400 4102
<< locali >>
rect 5946 4129 6214 4130
rect 4902 4085 6214 4129
rect 4902 4084 5991 4085
rect 4902 4022 4947 4084
rect 5417 4030 5462 4084
rect 5946 4020 5991 4084
rect 4721 3872 4819 3906
rect 4597 3613 4631 3727
rect 4721 3679 4755 3872
rect 4878 3679 4923 3748
rect 5459 3679 5504 3754
rect 5878 3679 5923 3752
rect 6169 3679 6214 4085
rect 6297 4062 6331 4221
rect 7179 4200 12383 4246
rect 7700 3996 7734 4200
rect 7870 4099 8756 4133
rect 7870 4043 7905 4099
rect 8722 4052 8756 4099
rect 9698 3970 9738 4200
rect 6324 3820 6454 3914
rect 3546 2141 3660 3206
rect 4685 3095 4791 3679
rect 4878 3634 6214 3679
rect 6297 3559 6331 3716
rect 5864 3525 6331 3559
rect 5864 3446 5898 3525
rect 6541 3401 6575 3748
rect 6982 3404 7230 3698
rect 8140 3408 8462 3752
rect 8733 3713 9617 3967
rect 3874 2420 4306 2576
rect 5176 2568 5608 2724
rect 5176 2246 5608 2402
rect 3876 2064 4308 2220
rect 4050 1796 5194 1912
rect 5864 1635 5898 1718
rect 6487 1635 6521 1753
rect 7185 1635 7219 1753
rect 7971 1635 8005 1755
rect 8753 1635 8787 1755
rect 9126 1635 9160 1718
rect 5864 1601 9160 1635
rect 9363 1512 9617 3713
rect 9698 3506 9732 3970
rect 10225 3925 10271 4200
rect 10766 3970 10800 4200
rect 10788 3802 11082 3936
rect 11467 3913 11513 4200
rect 11924 3954 11958 4200
rect 11762 3902 11945 3936
rect 11821 3868 11856 3902
rect 10148 3470 10406 3788
rect 11170 3784 11255 3818
rect 10766 3635 10800 3762
rect 10766 3601 10994 3635
rect 10960 3506 10994 3601
rect 11821 3603 11855 3843
rect 11924 3699 11958 3766
rect 11924 3665 12362 3699
rect 11821 3569 12259 3603
rect 11089 3434 11190 3468
rect 10986 3340 11082 3424
rect 12225 3409 12259 3569
rect 12328 3486 12362 3665
rect 10960 3211 10994 3298
rect 10540 3177 10994 3211
rect 10540 3046 10574 3177
rect 11450 3010 11574 3330
rect 9940 2628 10076 2826
rect 9774 1716 9910 1914
rect 10112 1734 10248 1932
rect 10406 1648 10506 1934
rect 10596 1684 10630 1712
rect 10596 1650 10680 1684
rect 10596 1649 10630 1650
rect 10736 1512 10794 1660
rect 10986 1512 11020 1632
rect 7500 1258 11345 1512
<< viali >>
rect 4685 2989 4791 3095
rect 3546 2027 3660 2141
<< metal1 >>
rect 8058 4020 8478 4344
rect 4310 3682 4362 3928
rect 6046 3866 6252 3918
rect 3015 3630 4362 3682
rect 4310 3588 4362 3630
rect 5961 3588 6007 3589
rect 6200 3588 6252 3866
rect 9504 3836 9822 3888
rect 9504 3588 9556 3836
rect 11318 3770 11420 3794
rect 11318 3662 11420 3668
rect 4310 3536 9556 3588
rect 5961 3366 6007 3536
rect 9496 3346 9844 3426
rect 9224 3316 9304 3322
rect 9496 3316 9576 3346
rect 4527 3252 5016 3316
rect 4483 3236 5016 3252
rect 5096 3236 5102 3316
rect 9304 3236 9576 3316
rect 4483 3041 4537 3236
rect 9224 3230 9304 3236
rect 9711 3127 9717 3229
rect 9819 3127 9825 3229
rect 3093 2987 4537 3041
rect 4673 3095 4803 3101
rect 4673 2989 4685 3095
rect 4791 2989 4803 3095
rect 4673 2983 4803 2989
rect 4685 2813 4791 2983
rect 9717 2825 9819 3127
rect 11029 2992 11350 3026
rect 3877 2707 4791 2813
rect 10264 2510 10464 2606
rect 10368 2170 10464 2510
rect 3534 2141 3672 2147
rect 3534 2027 3546 2141
rect 3660 2027 3672 2141
rect 5176 2036 5827 2106
rect 10368 2074 10800 2170
rect 3534 2021 3672 2027
rect 3546 1615 3660 2021
rect 5246 803 5360 1674
rect 5757 1518 5827 2036
rect 10704 1926 10800 2074
rect 5757 1447 8359 1518
rect 8288 781 8359 1447
<< via1 >>
rect 11318 3668 11420 3770
rect 5016 3236 5096 3316
rect 9224 3236 9304 3316
rect 9717 3127 9819 3229
<< metal2 >>
rect 11312 3668 11318 3770
rect 11420 3668 11426 3770
rect 5016 3316 5096 3322
rect 5096 3236 9224 3316
rect 9304 3236 9310 3316
rect 5016 3230 5096 3236
rect 9717 3229 9819 3235
rect 11318 3229 11420 3668
rect 9819 3127 11420 3229
rect 9717 3121 9819 3127
use M1  M1_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713519087
transform 0 1 11510 -1 0 3860
box -226 -484 226 484
use M2  M2_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713519243
transform 0 1 11714 -1 0 3392
box -226 -684 226 684
use M3  M3_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713519362
transform 0 -1 10848 1 0 2932
box -246 -344 246 344
use M3  M3_1
timestamp 1713519362
transform 0 1 11534 -1 0 2930
box -246 -344 246 344
use M7  M7_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713518916
transform 0 -1 10757 -1 0 1796
box -296 -299 296 299
use M9  M9_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713524830
transform 0 -1 10252 1 0 3866
box -236 -584 236 584
use M10  M10_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713518505
transform 0 -1 10346 -1 0 3402
box -236 -684 236 684
use M14  M14_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713520534
transform 0 1 5443 -1 0 3889
box -305 -919 305 1002
use M16  M16_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713520667
transform 0 -1 7512 -1 0 2582
box -996 -1684 996 1684
use M19  M19_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713520772
transform 0 -1 7086 -1 0 3832
box -296 -684 296 684
use M27  M27_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713522689
transform 0 1 8313 -1 0 3888
box -296 -479 296 479
use p7  p7_0
timestamp 1713528272
transform 1 0 12 0 1 1416
box -12 -1416 7768 2830
use Q2  Q2_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713441746
transform 1 0 2 0 1 -600
box 7780 600 9120 1940
use sky130_fd_pr__res_high_po_0p35_CMWQMJ  sky130_fd_pr__res_high_po_0p35_CMWQMJ_0
timestamp 0
transform 0 1 4742 -1 0 2403
box -533 -1032 533 1032
use sky130_fd_pr__res_high_po_0p35_K2NARC  sky130_fd_pr__res_high_po_0p35_K2NARC_0
timestamp 0
transform 1 0 10008 0 1 2278
box -450 -828 450 828
use sky130_fd_pr__res_high_po_0p35_N7UQCW  sky130_fd_pr__res_high_po_0p35_N7UQCW_0
timestamp 0
transform 0 1 4449 -1 0 1649
box -201 -1237 201 1237
<< end >>

magic
tech sky130B
magscale 1 2
timestamp 1713559273
<< metal4 >>
rect -2849 6239 2849 6280
rect -2849 161 2593 6239
rect 2829 161 2849 6239
rect -2849 120 2849 161
rect -2849 -161 2849 -120
rect -2849 -6239 2593 -161
rect 2829 -6239 2849 -161
rect -2849 -6280 2849 -6239
<< via4 >>
rect 2593 161 2829 6239
rect 2593 -6239 2829 -161
<< mimcap2 >>
rect -2769 6160 2231 6200
rect -2769 240 -2729 6160
rect 2191 240 2231 6160
rect -2769 200 2231 240
rect -2769 -240 2231 -200
rect -2769 -6160 -2729 -240
rect 2191 -6160 2231 -240
rect -2769 -6200 2231 -6160
<< mimcap2contact >>
rect -2729 240 2191 6160
rect -2729 -6160 2191 -240
<< metal5 >>
rect -429 6184 -109 6400
rect 2551 6239 2871 6400
rect -2753 6160 2215 6184
rect -2753 240 -2729 6160
rect 2191 240 2215 6160
rect -2753 216 2215 240
rect -429 -216 -109 216
rect 2551 161 2593 6239
rect 2829 161 2871 6239
rect 2551 -161 2871 161
rect -2753 -240 2215 -216
rect -2753 -6160 -2729 -240
rect 2191 -6160 2215 -240
rect -2753 -6184 2215 -6160
rect -429 -6400 -109 -6184
rect 2551 -6239 2593 -161
rect 2829 -6239 2871 -161
rect 2551 -6400 2871 -6239
<< properties >>
string FIXED_BBOX -2849 120 2311 6280
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 25 l 30 val 1.52k carea 2.00 cperi 0.19 nx 1 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

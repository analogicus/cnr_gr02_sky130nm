magic
tech sky130B
magscale 1 2
timestamp 1713559273
<< metal4 >>
rect -10447 6239 -3749 6280
rect -10447 161 -4005 6239
rect -3769 161 -3749 6239
rect -10447 120 -3749 161
rect -3349 6239 3349 6280
rect -3349 161 3093 6239
rect 3329 161 3349 6239
rect -3349 120 3349 161
rect 3749 6239 10447 6280
rect 3749 161 10191 6239
rect 10427 161 10447 6239
rect 3749 120 10447 161
rect -10447 -161 -3749 -120
rect -10447 -6239 -4005 -161
rect -3769 -6239 -3749 -161
rect -10447 -6280 -3749 -6239
rect -3349 -161 3349 -120
rect -3349 -6239 3093 -161
rect 3329 -6239 3349 -161
rect -3349 -6280 3349 -6239
rect 3749 -161 10447 -120
rect 3749 -6239 10191 -161
rect 10427 -6239 10447 -161
rect 3749 -6280 10447 -6239
<< via4 >>
rect -4005 161 -3769 6239
rect 3093 161 3329 6239
rect 10191 161 10427 6239
rect -4005 -6239 -3769 -161
rect 3093 -6239 3329 -161
rect 10191 -6239 10427 -161
<< mimcap2 >>
rect -10367 6160 -4367 6200
rect -10367 240 -10327 6160
rect -4407 240 -4367 6160
rect -10367 200 -4367 240
rect -3269 6160 2731 6200
rect -3269 240 -3229 6160
rect 2691 240 2731 6160
rect -3269 200 2731 240
rect 3829 6160 9829 6200
rect 3829 240 3869 6160
rect 9789 240 9829 6160
rect 3829 200 9829 240
rect -10367 -240 -4367 -200
rect -10367 -6160 -10327 -240
rect -4407 -6160 -4367 -240
rect -10367 -6200 -4367 -6160
rect -3269 -240 2731 -200
rect -3269 -6160 -3229 -240
rect 2691 -6160 2731 -240
rect -3269 -6200 2731 -6160
rect 3829 -240 9829 -200
rect 3829 -6160 3869 -240
rect 9789 -6160 9829 -240
rect 3829 -6200 9829 -6160
<< mimcap2contact >>
rect -10327 240 -4407 6160
rect -3229 240 2691 6160
rect 3869 240 9789 6160
rect -10327 -6160 -4407 -240
rect -3229 -6160 2691 -240
rect 3869 -6160 9789 -240
<< metal5 >>
rect -7527 6184 -7207 6400
rect -4047 6239 -3727 6400
rect -10351 6160 -4383 6184
rect -10351 240 -10327 6160
rect -4407 240 -4383 6160
rect -10351 216 -4383 240
rect -7527 -216 -7207 216
rect -4047 161 -4005 6239
rect -3769 161 -3727 6239
rect -429 6184 -109 6400
rect 3051 6239 3371 6400
rect -3253 6160 2715 6184
rect -3253 240 -3229 6160
rect 2691 240 2715 6160
rect -3253 216 2715 240
rect -4047 -161 -3727 161
rect -10351 -240 -4383 -216
rect -10351 -6160 -10327 -240
rect -4407 -6160 -4383 -240
rect -10351 -6184 -4383 -6160
rect -7527 -6400 -7207 -6184
rect -4047 -6239 -4005 -161
rect -3769 -6239 -3727 -161
rect -429 -216 -109 216
rect 3051 161 3093 6239
rect 3329 161 3371 6239
rect 6669 6184 6989 6400
rect 10149 6239 10469 6400
rect 3845 6160 9813 6184
rect 3845 240 3869 6160
rect 9789 240 9813 6160
rect 3845 216 9813 240
rect 3051 -161 3371 161
rect -3253 -240 2715 -216
rect -3253 -6160 -3229 -240
rect 2691 -6160 2715 -240
rect -3253 -6184 2715 -6160
rect -4047 -6400 -3727 -6239
rect -429 -6400 -109 -6184
rect 3051 -6239 3093 -161
rect 3329 -6239 3371 -161
rect 6669 -216 6989 216
rect 10149 161 10191 6239
rect 10427 161 10469 6239
rect 10149 -161 10469 161
rect 3845 -240 9813 -216
rect 3845 -6160 3869 -240
rect 9789 -6160 9813 -240
rect 3845 -6184 9813 -6160
rect 3051 -6400 3371 -6239
rect 6669 -6400 6989 -6184
rect 10149 -6239 10191 -161
rect 10427 -6239 10469 -161
rect 10149 -6400 10469 -6239
<< properties >>
string FIXED_BBOX 3749 120 9909 6280
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 3 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

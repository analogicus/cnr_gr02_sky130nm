magic
tech sky130B
magscale 1 2
timestamp 1713555407
<< nwell >>
rect 802 2054 1890 2286
<< locali >>
rect 1282 2784 1961 2830
rect 1282 2525 1328 2784
rect 1910 2566 1944 2784
rect 778 2428 858 2482
rect 1910 2285 1944 2358
rect 1809 2251 1944 2285
rect 1809 1947 1843 2251
<< metal1 >>
rect 1250 1940 1366 2382
rect 1799 1792 1851 2438
rect 1688 1740 1851 1792
use M9  M9_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713524830
transform 0 1 1396 -1 0 2462
box -236 -584 236 584
use p2  p2_0
timestamp 1713555407
transform 1 0 0 0 1 0
box 0 0 1878 2830


magic
tech sky130B
magscale 1 2
timestamp 1714173242
<< locali >>
rect 4608 5170 4992 5176
rect 4608 4856 4614 5170
rect -111 4798 4614 4856
rect 4986 4798 4992 5170
rect -111 4577 4992 4798
rect -111 1313 168 4577
rect 4608 4524 4992 4577
rect 247 4235 17012 4425
rect 4351 4200 5278 4235
rect 12852 3264 12982 3913
rect 16822 3204 17012 4235
rect 4685 3111 5279 3201
rect 4685 3095 5393 3111
rect 5173 3005 5393 3095
rect 12335 2871 12441 2877
rect 10931 2667 10997 2863
rect 11513 2669 11579 2855
rect 12335 2777 12341 2871
rect 12435 2777 12441 2871
rect 10931 2601 11392 2667
rect 11513 2603 12118 2669
rect 11326 1890 11392 2601
rect 12052 1888 12118 2603
rect 12335 2187 12441 2777
rect 12335 2081 12619 2187
rect 12513 2057 12619 2081
rect 12513 1951 12935 2057
rect 11006 1696 11112 1838
rect 11672 1730 11778 1872
rect 11320 1512 11416 1658
rect 11649 1512 11683 1633
rect 11752 1512 11786 1632
rect 12042 1512 12148 1666
rect 12304 1512 12338 1632
rect 11091 1258 12677 1512
rect 12423 152 12677 1258
rect 12422 -40 12946 152
<< viali >>
rect 4614 4798 4986 5170
rect 5393 3005 5499 3111
rect 12341 2777 12435 2871
<< metal1 >>
rect 4132 5176 4516 5182
rect 4516 5170 4998 5176
rect 4516 4798 4614 5170
rect 4986 4798 4998 5170
rect 4516 4792 4998 4798
rect 7414 5108 7734 5114
rect 4132 4786 4516 4792
rect 7414 4620 7734 4788
rect 7414 4340 8488 4620
rect 7414 4300 12676 4340
rect 8428 4236 12676 4300
rect 5387 3111 5505 3123
rect 5387 3005 5393 3111
rect 5499 3005 5603 3111
rect 5709 3005 5715 3111
rect 12335 3045 12441 3051
rect 5387 2993 5505 3005
rect 12335 2871 12441 2939
rect 12335 2777 12341 2871
rect 12435 2777 12441 2871
rect 12335 2765 12441 2777
rect 12572 2592 12676 4236
rect 12572 2488 12926 2592
rect 11570 1750 11872 1800
<< via1 >>
rect 4132 4792 4516 5176
rect 7414 4788 7734 5108
rect 5603 3005 5709 3111
rect 12335 2939 12441 3045
<< metal2 >>
rect 3671 5176 4045 5180
rect 3666 5171 4132 5176
rect 3666 4797 3671 5171
rect 4045 4797 4132 5171
rect 3666 4792 4132 4797
rect 4516 4792 4522 5176
rect 7859 5108 8169 5112
rect 3671 4788 4045 4792
rect 7408 4788 7414 5108
rect 7734 5103 8174 5108
rect 7734 4793 7859 5103
rect 8169 4793 8174 5103
rect 7734 4788 8174 4793
rect 7859 4784 8169 4788
rect 5603 3111 5709 3117
rect 5709 3045 9645 3111
rect 5709 3005 12335 3045
rect 5603 2999 5709 3005
rect 9539 2939 12335 3005
rect 12441 2939 12447 3045
<< via2 >>
rect 3671 4797 4045 5171
rect 7859 4793 8169 5103
<< metal3 >>
rect 3098 5175 4050 5176
rect 3093 4793 3099 5175
rect 3481 5171 4050 5175
rect 3481 4797 3671 5171
rect 4045 4797 4050 5171
rect 8311 5108 8629 5113
rect 3481 4793 4050 4797
rect 3098 4792 4050 4793
rect 7854 5107 8630 5108
rect 7854 5103 8311 5107
rect 7854 4793 7859 5103
rect 8169 4793 8311 5103
rect 7854 4789 8311 4793
rect 8629 4789 8630 5107
rect 7854 4788 8630 4789
rect 8311 4783 8629 4788
<< via3 >>
rect 3099 4793 3481 5175
rect 8311 4789 8629 5107
<< metal4 >>
rect 1518 18720 8158 19012
rect 1518 17612 1810 18720
rect 1446 16880 1810 17612
rect 1446 9134 1738 16880
rect 7866 14310 8158 18720
rect 7866 14018 16356 14310
rect 16064 9134 16356 14018
rect 1446 8842 16356 9134
rect 3098 5175 3482 5572
rect 3098 4793 3099 5175
rect 3481 4793 3482 5175
rect 3098 4792 3482 4793
rect 8310 5107 9242 5108
rect 8310 4789 8311 5107
rect 8629 5084 9242 5107
rect 8629 4812 8946 5084
rect 9218 4812 9242 5084
rect 8629 4789 9242 4812
rect 8310 4788 9242 4789
<< via4 >>
rect 8946 4812 9218 5084
<< metal5 >>
rect 3940 19584 4260 19592
rect 3940 19264 7658 19584
rect 3940 8208 4260 19264
rect 7338 15202 7658 19264
rect 7338 14988 16802 15202
rect 7344 14882 16802 14988
rect 16482 8208 16802 14882
rect 3932 7888 16802 8208
rect 8922 5084 9242 5506
rect 8922 4812 8946 5084
rect 9218 4812 9242 5084
rect 8922 4788 9242 4812
use COMP  COMP_0
timestamp 1713519326
transform 0 1 15962 -1 0 -2716
box -6200 -3190 -2588 1050
use M6  M6_0
timestamp 1713519460
transform 0 1 11390 -1 0 1777
box -276 -329 276 329
use M6  M6_1
timestamp 1713519460
transform 0 -1 12045 -1 0 1776
box -276 -329 276 329
use P16  P16_0
timestamp 1713561060
transform 1 0 0 0 1 0
box 0 0 12400 4344
use sky130_fd_pr__cap_mim_m3_2_L4ZKLG  sky130_fd_pr__cap_mim_m3_2_L4ZKLG_0
timestamp 1713559273
transform 1 0 6890 0 1 11594
box -6898 -6400 6920 6400
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_0
timestamp 1713559273
transform 1 0 3371 0 1 21563
box -3349 -3081 3371 3081
use sky130_fd_pr__cap_mim_m3_2_M9XTT6  sky130_fd_pr__cap_mim_m3_2_M9XTT6_0
timestamp 1713559273
transform 1 0 8828 0 1 21561
box -1778 -3081 1800 3081
use sky130_fd_pr__cap_mim_m3_2_SJC7NT  sky130_fd_pr__cap_mim_m3_2_SJC7NT_0
timestamp 1713559273
transform 1 0 16911 0 1 11628
box -2849 -6400 2871 6400
<< labels >>
flabel locali 380 4294 772 4388 0 FreeSans 800 0 0 0 VDD_1V8
port 0 nsew
flabel locali 118 1374 510 1468 0 FreeSans 800 0 0 0 VSS
port 1 nsew
flabel locali 12866 3508 12962 3880 0 FreeSans 800 0 0 0 VO
port 2 nsew
flabel locali 8628 3818 8646 3954 0 FreeSans 400 0 0 0 rst
port 3 nsew
flabel locali 11336 2230 11378 2448 0 FreeSans 400 0 0 0 LPO
port 4 nsew
flabel locali 770 1960 790 2186 0 FreeSans 400 0 0 0 LPI
port 6 nsew
<< end >>

magic
tech sky130B
timestamp 1713476524
<< pwell >>
rect -100 -586 100 586
<< psubdiff >>
rect -82 520 -65 551
rect -82 -551 -65 -520
<< psubdiffcont >>
rect -82 -520 -65 520
<< xpolycontact >>
rect -17 287 17 503
rect -17 -503 17 -287
<< ppolyres >>
rect -17 -287 17 287
<< locali >>
rect -82 520 -65 551
rect -82 -551 -65 -520
<< viali >>
rect -9 295 9 494
rect -9 -494 9 -295
<< metal1 >>
rect -12 494 12 500
rect -12 295 -9 494
rect 9 295 12 494
rect -12 289 12 295
rect -12 -295 12 -289
rect -12 -494 -9 -295
rect 9 -494 12 -295
rect -12 -500 12 -494
<< properties >>
string FIXED_BBOX -74 -559 74 559
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.35 l 5.9 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 6.504k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

magic
tech sky130B
magscale 1 2
timestamp 1713559273
<< metal4 >>
rect -6898 6239 -200 6280
rect -6898 161 -456 6239
rect -220 161 -200 6239
rect -6898 120 -200 161
rect 200 6239 6898 6280
rect 200 161 6642 6239
rect 6878 161 6898 6239
rect 200 120 6898 161
rect -6898 -161 -200 -120
rect -6898 -6239 -456 -161
rect -220 -6239 -200 -161
rect -6898 -6280 -200 -6239
rect 200 -161 6898 -120
rect 200 -6239 6642 -161
rect 6878 -6239 6898 -161
rect 200 -6280 6898 -6239
<< via4 >>
rect -456 161 -220 6239
rect 6642 161 6878 6239
rect -456 -6239 -220 -161
rect 6642 -6239 6878 -161
<< mimcap2 >>
rect -6818 6160 -818 6200
rect -6818 240 -6778 6160
rect -858 240 -818 6160
rect -6818 200 -818 240
rect 280 6160 6280 6200
rect 280 240 320 6160
rect 6240 240 6280 6160
rect 280 200 6280 240
rect -6818 -240 -818 -200
rect -6818 -6160 -6778 -240
rect -858 -6160 -818 -240
rect -6818 -6200 -818 -6160
rect 280 -240 6280 -200
rect 280 -6160 320 -240
rect 6240 -6160 6280 -240
rect 280 -6200 6280 -6160
<< mimcap2contact >>
rect -6778 240 -858 6160
rect 320 240 6240 6160
rect -6778 -6160 -858 -240
rect 320 -6160 6240 -240
<< metal5 >>
rect -3978 6184 -3658 6400
rect -498 6239 -178 6400
rect -6802 6160 -834 6184
rect -6802 240 -6778 6160
rect -858 240 -834 6160
rect -6802 216 -834 240
rect -3978 -216 -3658 216
rect -498 161 -456 6239
rect -220 161 -178 6239
rect 3120 6184 3440 6400
rect 6600 6239 6920 6400
rect 296 6160 6264 6184
rect 296 240 320 6160
rect 6240 240 6264 6160
rect 296 216 6264 240
rect -498 -161 -178 161
rect -6802 -240 -834 -216
rect -6802 -6160 -6778 -240
rect -858 -6160 -834 -240
rect -6802 -6184 -834 -6160
rect -3978 -6400 -3658 -6184
rect -498 -6239 -456 -161
rect -220 -6239 -178 -161
rect 3120 -216 3440 216
rect 6600 161 6642 6239
rect 6878 161 6920 6239
rect 6600 -161 6920 161
rect 296 -240 6264 -216
rect 296 -6160 320 -240
rect 6240 -6160 6264 -240
rect 296 -6184 6264 -6160
rect -498 -6400 -178 -6239
rect 3120 -6400 3440 -6184
rect 6600 -6239 6642 -161
rect 6878 -6239 6920 -161
rect 6600 -6400 6920 -6239
<< properties >>
string FIXED_BBOX 200 120 6360 6280
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

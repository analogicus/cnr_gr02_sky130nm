magic
tech sky130B
magscale 1 2
timestamp 1713258660
<< error_s >>
rect 36258 5434 36482 5436
rect 19670 2376 19704 2430
rect 10382 1941 10454 1947
rect 10520 1941 10592 1947
rect 7807 626 7809 1914
rect 10382 1907 10394 1941
rect 10520 1907 10532 1941
rect 10382 1901 10454 1907
rect 10520 1901 10592 1907
rect 10691 1628 10792 1882
rect 9050 1385 9095 1403
rect 9050 1349 9222 1385
rect 9068 753 9222 1349
rect 9607 1315 9642 1349
rect 9608 1296 9642 1315
rect 9268 1247 9340 1253
rect 9406 1247 9478 1253
rect 9268 1213 9280 1247
rect 9406 1213 9418 1247
rect 9268 1207 9340 1213
rect 9406 1207 9478 1213
rect 9068 626 9138 753
rect 9268 719 9340 725
rect 9406 719 9478 725
rect 9268 685 9280 719
rect 9406 685 9418 719
rect 9268 679 9340 685
rect 9406 679 9478 685
rect 9068 600 9129 626
rect 9104 592 9129 600
rect 9627 583 9642 1296
rect 9661 1262 9696 1296
rect 9661 583 9695 1262
rect 9825 1194 9897 1200
rect 9963 1194 10035 1200
rect 9825 1160 9837 1194
rect 9963 1160 9975 1194
rect 9825 1154 9897 1160
rect 9963 1154 10035 1160
rect 9825 666 9897 672
rect 9963 666 10035 672
rect 9825 632 9837 666
rect 9963 632 9975 666
rect 9825 626 9897 632
rect 9963 626 10035 632
rect 9661 549 9676 583
rect 10184 530 10199 1296
rect 10218 530 10252 1350
rect 10382 613 10454 619
rect 10520 613 10592 619
rect 10382 579 10394 613
rect 10520 579 10532 613
rect 10945 594 11046 1628
rect 12079 594 12233 1882
rect 15659 1037 15693 1091
rect 10382 573 10454 579
rect 10520 573 10592 579
rect 10218 496 10233 530
rect 12079 467 12149 594
rect 12079 441 12140 467
rect 12115 433 12140 441
rect 15678 424 15693 1037
rect 15712 1003 15747 1037
rect 15712 424 15746 1003
rect 15873 935 15931 941
rect 15991 935 16049 941
rect 15873 901 15885 935
rect 15991 901 16003 935
rect 15873 895 15931 901
rect 15991 895 16049 901
rect 15873 507 15931 513
rect 15991 507 16049 513
rect 15873 473 15885 507
rect 15991 473 16003 507
rect 15873 467 15931 473
rect 15991 467 16049 473
rect 15712 390 15727 424
rect 16195 371 16210 1037
rect 16229 371 16263 1088
rect 16390 1082 16448 1088
rect 16508 1082 16566 1088
rect 16390 1048 16402 1082
rect 16508 1048 16520 1082
rect 16390 1042 16448 1048
rect 16508 1042 16566 1048
rect 16693 791 16727 845
rect 16390 454 16448 460
rect 16508 454 16566 460
rect 16390 420 16402 454
rect 16508 420 16520 454
rect 16390 414 16448 420
rect 16508 414 16566 420
rect 16229 337 16244 371
rect 16712 318 16727 791
rect 16746 757 16781 791
rect 17289 757 17324 791
rect 16746 318 16780 757
rect 17290 738 17324 757
rect 16746 284 16761 318
rect 17309 265 17324 738
rect 17343 704 17378 738
rect 17886 704 17921 711
rect 17343 265 17377 704
rect 17887 693 17921 704
rect 17887 657 17957 693
rect 17904 623 17975 657
rect 18603 623 18638 657
rect 17343 231 17358 265
rect 17904 212 17974 623
rect 18604 604 18638 623
rect 17904 176 17957 212
rect 18623 159 18638 604
rect 18657 570 18692 604
rect 18657 159 18691 570
rect 18657 125 18672 159
rect 19340 106 19355 604
rect 19374 106 19408 658
rect 19374 72 19389 106
rect 19689 53 19704 2376
rect 19723 2342 19758 2376
rect 19723 53 19757 2342
rect 23372 567 23407 601
rect 23875 567 23910 601
rect 20019 415 20053 469
rect 19723 19 19738 53
rect 20038 0 20053 415
rect 20072 381 20107 415
rect 20072 0 20106 381
rect 20072 -34 20087 0
rect 20835 -53 20850 415
rect 20869 -53 20903 469
rect 22979 452 23051 458
rect 23117 452 23189 458
rect 21165 389 21199 443
rect 22815 425 22849 443
rect 20869 -87 20884 -53
rect 21184 -106 21199 389
rect 21218 355 21253 389
rect 21218 -106 21252 355
rect 21218 -140 21233 -106
rect 22779 -159 22849 425
rect 22979 418 22991 452
rect 23117 418 23129 452
rect 22979 412 23051 418
rect 23117 412 23189 418
rect 22979 -76 23051 -70
rect 23117 -76 23189 -70
rect 22979 -110 22991 -76
rect 23117 -110 23129 -76
rect 22979 -116 23051 -110
rect 23117 -116 23189 -110
rect 22779 -195 22832 -159
rect 23338 -212 23353 554
rect 23372 -212 23406 567
rect 23876 548 23910 567
rect 23536 499 23608 505
rect 23674 499 23746 505
rect 23536 465 23548 499
rect 23674 465 23686 499
rect 23536 459 23608 465
rect 23674 459 23746 465
rect 23536 -129 23608 -123
rect 23674 -129 23746 -123
rect 23536 -163 23548 -129
rect 23674 -163 23686 -129
rect 23536 -169 23608 -163
rect 23674 -169 23746 -163
rect 23372 -246 23387 -212
rect 23895 -265 23910 548
rect 23929 514 23964 548
rect 24432 514 24467 548
rect 23929 -265 23963 514
rect 24433 495 24467 514
rect 24093 446 24165 452
rect 24231 446 24303 452
rect 24093 412 24105 446
rect 24231 412 24243 446
rect 24093 406 24165 412
rect 24231 406 24303 412
rect 24093 -182 24165 -176
rect 24231 -182 24303 -176
rect 24093 -216 24105 -182
rect 24231 -216 24243 -182
rect 24093 -222 24165 -216
rect 24231 -222 24303 -216
rect 23929 -299 23944 -265
rect 24452 -318 24467 495
rect 24486 461 24521 495
rect 24486 -318 24520 461
rect 24650 393 24722 399
rect 24788 393 24860 399
rect 24650 359 24662 393
rect 24788 359 24800 393
rect 24650 353 24722 359
rect 24788 353 24860 359
rect 28391 196 28426 230
rect 28894 196 28929 230
rect 27834 154 27869 172
rect 27798 149 27869 154
rect 24990 42 25024 96
rect 27037 84 27072 95
rect 25804 42 25857 77
rect 24650 -235 24722 -229
rect 24788 -235 24860 -229
rect 24650 -269 24662 -235
rect 24788 -269 24800 -235
rect 24650 -275 24722 -269
rect 24788 -275 24860 -269
rect 24486 -352 24501 -318
rect 25009 -371 25024 42
rect 25043 8 25078 42
rect 25786 41 25857 42
rect 25043 -371 25077 8
rect 25804 7 25875 41
rect 25043 -405 25058 -371
rect 25804 -424 25874 7
rect 25804 -460 25857 -424
rect 27003 -477 27018 41
rect 27037 -477 27071 84
rect 27037 -511 27052 -477
rect 27798 -530 27868 149
rect 27998 81 28070 87
rect 28136 81 28208 87
rect 27998 47 28010 81
rect 28136 47 28148 81
rect 27998 41 28070 47
rect 28136 41 28208 47
rect 27998 -447 28070 -441
rect 28136 -447 28208 -441
rect 27998 -481 28010 -447
rect 28136 -481 28148 -447
rect 27998 -487 28070 -481
rect 28136 -487 28208 -481
rect 27798 -566 27851 -530
rect 28357 -583 28372 183
rect 28391 -583 28425 196
rect 28895 177 28929 196
rect 28555 128 28627 134
rect 28693 128 28765 134
rect 28555 94 28567 128
rect 28693 94 28705 128
rect 28555 88 28627 94
rect 28693 88 28765 94
rect 28555 -500 28627 -494
rect 28693 -500 28765 -494
rect 28555 -534 28567 -500
rect 28693 -534 28705 -500
rect 28555 -540 28627 -534
rect 28693 -540 28765 -534
rect 28391 -617 28406 -583
rect 28914 -636 28929 177
rect 28948 143 28983 177
rect 28948 -636 28982 143
rect 28948 -670 28963 -636
rect 36258 -726 36540 5434
rect 42978 5433 43202 5435
rect 36578 -630 36802 5338
rect 42978 -727 43260 5433
rect 49698 5432 49922 5434
rect 43298 -631 43522 5337
rect 49698 -728 49980 5432
rect 56418 5431 56642 5433
rect 50018 -632 50242 5336
rect 56418 -729 56700 5431
rect 63138 5430 63362 5432
rect 56738 -633 56962 5335
rect 63138 -730 63420 5430
rect 63458 -634 63682 5334
rect 69858 1429 70082 1653
rect 72802 1430 72860 1509
rect 69858 -731 70140 1429
rect 70178 -635 70402 1333
rect 72578 -732 72860 1430
rect 72898 -636 73122 1750
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__cap_mim_m3_2_3HBNLG  XC1
timestamp 1713258222
transform 1 0 33111 0 1 2355
box -3349 -3081 3371 3081
use sky130_fd_pr__cap_mim_m3_2_3HBNLG  XC2
timestamp 1713258222
transform 1 0 39831 0 1 2354
box -3349 -3081 3371 3081
use sky130_fd_pr__cap_mim_m3_2_3HBNLG  XC3
timestamp 1713258222
transform 1 0 46551 0 1 2353
box -3349 -3081 3371 3081
use sky130_fd_pr__cap_mim_m3_2_3HBNLG  XC4
timestamp 1713258222
transform 1 0 53271 0 1 2352
box -3349 -3081 3371 3081
use sky130_fd_pr__cap_mim_m3_2_3HBNLG  XC5
timestamp 1713258222
transform 1 0 59991 0 1 2351
box -3349 -3081 3371 3081
use sky130_fd_pr__cap_mim_m3_2_3HBNLG  XC6
timestamp 1713258222
transform 1 0 66711 0 1 2350
box -3349 -3081 3371 3081
use sky130_fd_pr__cap_mim_m3_2_4PHTN9  XC7
timestamp 1713258222
transform 1 0 71431 0 1 349
box -1349 -1081 1371 1081
use sky130_fd_pr__cap_mim_m3_2_3HBNLG  XC8
timestamp 1713258222
transform 1 0 76151 0 1 2348
box -3349 -3081 3371 3081
use sky130_fd_pr__pfet_01v8_JMC8WZ  XM1
timestamp 1713258222
transform 1 0 15961 0 1 704
box -285 -369 285 369
use sky130_fd_pr__pfet_01v8_JMP7WZ  XM2
timestamp 1713258222
transform 1 0 16478 0 1 751
box -285 -469 285 469
use sky130_fd_pr__pfet_01v8_XG4SY6  XM3
timestamp 1713258222
transform 1 0 17035 0 1 528
box -325 -299 325 299
use sky130_fd_pr__pfet_01v8_XG4SY6  XM4
timestamp 1713258222
transform 1 0 17632 0 1 475
box -325 -299 325 299
use sky130_fd_pr__nfet_01v8_U7AL37  XM5
timestamp 1713258222
transform 1 0 18289 0 1 408
box -385 -285 385 285
use sky130_fd_pr__nfet_01v8_U7AL37  XM6
timestamp 1713258222
transform 1 0 19006 0 1 355
box -385 -285 385 285
use sky130_fd_pr__nfet_01v8_ZYANF2  XM7
timestamp 1713258222
transform 1 0 20461 0 1 181
box -425 -270 425 270
use sky130_fd_pr__nfet_01v8_RFVHWA  XM8
timestamp 1713258222
transform 1 0 22007 0 1 115
box -825 -310 825 310
use sky130_fd_pr__pfet_01v8_XPP79A  XM9
timestamp 1713258222
transform 1 0 23084 0 1 171
box -305 -419 305 419
use sky130_fd_pr__pfet_01v8_TMP79A  XM10
timestamp 1713258222
transform 1 0 23641 0 1 168
box -305 -469 305 469
use sky130_fd_pr__pfet_01v8_TMP79A  XM11
timestamp 1713258222
transform 1 0 24198 0 1 115
box -305 -469 305 469
use sky130_fd_pr__pfet_01v8_XPP79A  XM12
timestamp 1713258222
transform 1 0 9373 0 1 966
box -305 -419 305 419
use sky130_fd_pr__pfet_01v8_XPP79A  XM13
timestamp 1713258222
transform 1 0 9930 0 1 913
box -305 -419 305 419
use sky130_fd_pr__pfet_01v8_XPB89A  XM14
timestamp 1713258222
transform 1 0 10487 0 1 1260
box -305 -819 305 819
use sky130_fd_pr__pfet_01v8_XPP79A  XM15
timestamp 1713258222
transform 1 0 28103 0 1 -200
box -305 -419 305 419
use sky130_fd_pr__pfet_01v8_CQBZVD  XM16
timestamp 1713258222
transform 1 0 13904 0 1 1357
box -1825 -969 1825 969
use sky130_fd_pr__pfet_01v8_TMP79A  XM17
timestamp 1713258222
transform 1 0 24755 0 1 62
box -305 -469 305 469
use sky130_fd_pr__pfet_01v8_TMP79A  XM18
timestamp 1713258222
transform 1 0 28660 0 1 -203
box -305 -469 305 469
use sky130_fd_pr__pfet_01v8_FQU9VM  XM19
timestamp 1713258222
transform 1 0 29337 0 1 -256
box -425 -469 425 469
use sky130_fd_pr__nfet_01v8_QGMQ49  XM20
timestamp 1713258222
transform 1 0 27426 0 1 -206
box -425 -360 425 360
use sky130_fd_pr__pfet_01v8_FQE7VM  XM21
timestamp 1713258222
transform 1 0 25432 0 1 -191
box -425 -269 425 269
use sky130_fd_pr__nfet_01v8_UTAWZB  XM22
timestamp 1713258222
transform 1 0 26429 0 1 -218
box -625 -295 625 295
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ1 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1705202102
transform 1 0 7781 0 1 600
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ2
array 0 5 1288 0 0 1288
timestamp 1705202102
transform 1 0 1 0 1 600
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ3
timestamp 1705202102
transform 1 0 10792 0 1 441
box 0 0 1340 1340
use sky130_fd_pr__res_high_po_0p35_WA83VQ  XR1
timestamp 1713258222
transform 1 0 19888 0 1 1188
box -201 -1224 201 1224
use sky130_fd_pr__res_high_po_0p35_WMUZZM  XR2
timestamp 1713258222
transform 1 0 19539 0 1 3281
box -201 -3264 201 3264
use sky130_fd_pr__res_high_po_0p35_HTJVTY  XR3
timestamp 1713258222
transform 1 0 21034 0 1 1761
box -201 -1903 201 1903
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD_1V8
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 rst
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VO
port 3 nsew
<< end >>

*----------------------------------------------------------------
* Include
*----------------------------------------------------------------

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TEMP=40 GMIN=1e-15 reltol=1e-6 abstol=1e-6 keepopinfo noopiter gminsteps=5

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p


*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD  0  dc 1.8
Vrst reset 0 pwl 0 1.8 10u 1.8 10.1u 0
Vop vop 0 pwl 0 1.8 20u 1.8 20.1u 0

Rd0 d0 VSS 1e6
Rd1 d1 VSS 1e6

adut [ clk reset vop ] [ rst d0 d1 d2 d3 d4 d5 d6 d7 d8 d9 d10 d11 d12 d13 d14 d15 ] null dut
.model dut d_cosim simulation="../../verilog/temp_to_digital.so"

 
.control

tran 100n 200u

save all
write
.endc
.end

magic
tech sky130B
timestamp 1715274076
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ2 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1698934549
transform 1 0 3890 0 1 300
box 0 0 670 670
<< end >>

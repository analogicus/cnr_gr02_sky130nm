magic
tech sky130B
magscale 1 2
timestamp 1715274076
<< error_p >>
rect -3762 -2376 -3731 -2272
rect -5023 -2431 -4961 -2403
rect -5013 -2484 -4966 -2437
rect -3524 -2791 -3477 -2744
<< locali >>
rect -6110 910 -4580 1050
rect -6110 830 -5920 910
rect -4770 830 -4580 910
rect -4540 870 -4250 1050
rect -4210 910 -2680 1050
rect -5960 440 -5680 670
rect -6000 -190 -5680 40
rect -5024 28 -4960 410
rect -5250 -102 -4986 -26
rect -4425 -44 -4354 870
rect -4210 830 -4020 910
rect -2870 830 -2680 910
rect -4120 410 -3800 640
rect -3365 493 -2927 559
rect -4426 -104 -4420 -44
rect -4360 -104 -4354 -44
rect -4426 -110 -4354 -104
rect -4120 -190 -3800 40
rect -3540 -106 -3536 -42
rect -3464 -106 -3058 -42
rect -6010 -800 -5690 -570
rect -5450 -710 -5446 -640
rect -5374 -710 -5370 -640
rect -5155 -689 -4970 -620
rect -6030 -1400 -5684 -1170
rect -5155 -1209 -5086 -689
rect -4100 -800 -3780 -570
rect -3124 -712 -3059 -203
rect -5278 -1278 -5086 -1209
rect -4100 -1400 -3780 -1170
rect -2993 -1247 -2927 493
rect -3123 -1313 -2927 -1247
rect -4525 -1691 -3179 -1685
rect -4525 -1749 -4519 -1691
rect -4461 -1749 -3179 -1691
rect -4525 -1755 -3179 -1749
rect -6030 -1990 -5684 -1760
rect -5264 -1866 -4982 -1801
rect -3958 -1846 -3894 -1840
rect -3958 -1898 -3952 -1846
rect -3900 -1898 -3894 -1846
rect -6030 -2590 -5684 -2360
rect -5463 -2450 -5109 -2387
rect -5023 -2431 -4961 -2005
rect -3958 -2138 -3894 -1898
rect -3958 -2202 -3762 -2138
rect -3245 -2143 -3183 -1755
rect -2866 -2051 -2677 -1350
rect -3826 -2306 -3762 -2202
rect -3641 -2205 -3183 -2143
rect -3765 -2376 -3762 -2306
rect -5172 -2786 -5109 -2450
rect -3826 -2606 -3762 -2376
rect -3118 -2469 -3065 -2309
rect -3246 -2522 -3065 -2469
rect -5861 -2848 -5108 -2786
rect -4392 -2848 -4329 -2672
rect -5861 -2849 -4329 -2848
rect -5861 -2980 -5798 -2849
rect -5172 -2911 -4329 -2849
rect -6110 -3110 -5600 -2980
rect -5460 -3039 -4950 -2980
rect -5460 -3080 -5247 -3039
rect -5206 -3080 -4950 -3039
rect -5460 -3110 -4950 -3080
rect -4840 -3034 -4330 -2980
rect -4840 -3083 -4684 -3034
rect -4635 -3083 -4330 -3034
rect -4840 -3110 -4330 -3083
rect -3246 -3164 -3193 -2522
rect -3122 -3029 -3061 -2905
rect -4296 -3171 -3193 -3164
rect -4296 -3212 -4291 -3171
rect -4250 -3200 -3193 -3171
rect -4250 -3212 -3194 -3200
rect -4296 -3217 -3194 -3212
<< viali >>
rect -5441 489 -5374 556
rect -5440 -110 -5380 -50
rect -3540 493 -3481 552
rect -4420 -104 -4360 -44
rect -3536 -110 -3464 -38
rect -5446 -710 -5374 -638
rect -3540 -686 -3476 -622
rect -5434 -1272 -5382 -1220
rect -5023 -1283 -4965 -1225
rect -3535 -1270 -3484 -1219
rect -4519 -1749 -4461 -1691
rect -5434 -1860 -5382 -1808
rect -3952 -1898 -3900 -1846
rect -5013 -2484 -4966 -2437
rect -4392 -2672 -4329 -2609
rect -3524 -2791 -3477 -2744
rect -5247 -3080 -5206 -3039
rect -4684 -3083 -4635 -3034
rect -3122 -3090 -3061 -3029
rect -4291 -3212 -4250 -3171
<< metal1 >>
rect -5447 558 -5368 568
rect -5447 556 -3469 558
rect -5447 489 -5441 556
rect -5374 552 -3469 556
rect -5374 493 -3540 552
rect -3481 493 -3469 552
rect -5374 489 -3469 493
rect -5447 487 -3469 489
rect -5447 477 -5368 487
rect -4426 -38 -4354 -32
rect -3542 -38 -3458 -26
rect -5446 -50 -5374 -38
rect -5446 -110 -5440 -50
rect -5380 -110 -5374 -50
rect -5446 -340 -5374 -110
rect -4426 -44 -3536 -38
rect -4426 -104 -4420 -44
rect -4360 -104 -3536 -44
rect -4426 -110 -3536 -104
rect -3464 -110 -3458 -38
rect -4426 -116 -4354 -110
rect -3542 -122 -3458 -110
rect -5450 -410 -4820 -340
rect -5446 -632 -5374 -410
rect -5458 -638 -5362 -632
rect -5458 -710 -5446 -638
rect -5374 -710 -5362 -638
rect -5458 -716 -5362 -710
rect -5440 -1220 -5376 -1208
rect -4890 -1219 -4820 -410
rect -3546 -622 -3470 -610
rect -5440 -1272 -5434 -1220
rect -5382 -1272 -5376 -1220
rect -5440 -1808 -5376 -1272
rect -5035 -1225 -4820 -1219
rect -5035 -1283 -5023 -1225
rect -4965 -1283 -4820 -1225
rect -5035 -1289 -4820 -1283
rect -4890 -1685 -4820 -1289
rect -4392 -686 -3540 -622
rect -3476 -686 -3470 -622
rect -4890 -1691 -4449 -1685
rect -4890 -1749 -4519 -1691
rect -4461 -1749 -4449 -1691
rect -4890 -1755 -4449 -1749
rect -5440 -1860 -5434 -1808
rect -5382 -1860 -5376 -1808
rect -5440 -1872 -5376 -1860
rect -4392 -1840 -4328 -686
rect -3546 -698 -3470 -686
rect -3547 -1219 -3179 -1213
rect -3547 -1270 -3535 -1219
rect -3484 -1270 -3179 -1219
rect -3547 -1276 -3179 -1270
rect -3958 -1840 -3894 -1834
rect -4392 -1846 -3894 -1840
rect -4392 -1898 -3952 -1846
rect -3900 -1898 -3894 -1846
rect -4392 -1904 -3894 -1898
rect -3958 -1910 -3894 -1904
rect -3242 -1959 -3179 -1276
rect -4391 -2022 -3179 -1959
rect -5019 -2437 -4960 -2425
rect -5019 -2484 -5013 -2437
rect -4966 -2484 -4960 -2437
rect -5019 -2738 -4960 -2484
rect -4391 -2603 -4328 -2022
rect -4404 -2609 -4317 -2603
rect -4404 -2672 -4392 -2609
rect -4329 -2672 -4317 -2609
rect -4404 -2678 -4317 -2672
rect -5019 -2744 -3465 -2738
rect -5019 -2791 -3524 -2744
rect -3477 -2791 -3465 -2744
rect -5019 -2797 -3465 -2791
rect -5253 -2939 -5200 -2916
rect -5253 -2992 -4864 -2939
rect -5253 -3039 -5200 -2992
rect -5253 -3080 -5247 -3039
rect -5206 -3080 -5200 -3039
rect -5253 -3092 -5200 -3080
rect -4917 -3165 -4864 -2992
rect -3134 -3028 -3049 -3023
rect -4696 -3029 -3049 -3028
rect -4696 -3034 -3122 -3029
rect -4696 -3083 -4684 -3034
rect -4635 -3083 -3122 -3034
rect -4696 -3089 -3122 -3083
rect -3134 -3090 -3122 -3089
rect -3061 -3090 -3049 -3029
rect -3134 -3096 -3049 -3090
rect -4917 -3171 -4238 -3165
rect -4917 -3212 -4291 -3171
rect -4250 -3212 -4238 -3171
rect -4917 -3218 -4238 -3212
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1712008800
transform 1 0 -4116 0 1 224
box -184 -124 1528 718
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_1
timestamp 1712008800
transform 1 0 -4116 0 1 -366
box -184 -124 1528 718
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_2
timestamp 1712008800
transform 1 0 -4116 0 1 -3066
box -184 -124 1528 718
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_3
timestamp 1712008800
transform 1 0 -4116 0 1 -956
box -184 -124 1528 718
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_4
timestamp 1712008800
transform 1 0 -4116 0 1 -2476
box -184 -124 1528 718
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_5
timestamp 1712008800
transform 1 0 -4116 0 1 -1546
box -184 -124 1528 718
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1712008800
transform 1 0 -6016 0 1 224
box -184 -124 1528 718
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_1
timestamp 1712008800
transform 1 0 -6016 0 1 -366
box -184 -124 1528 718
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_2
timestamp 1712008800
transform 1 0 -6016 0 1 -956
box -184 -124 1528 718
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_3
timestamp 1712008800
transform 1 0 -6016 0 1 -1546
box -184 -124 1528 718
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_4
timestamp 1712008800
transform 1 0 -6016 0 1 -2136
box -184 -124 1528 718
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_5
timestamp 1712008800
transform 1 0 -6016 0 1 -2726
box -184 -124 1528 718
<< labels >>
flabel locali -5670 930 -5000 1030 0 FreeSans 400 0 0 0 VDD
port 2 nsew
flabel locali -3850 920 -3030 1030 0 FreeSans 400 0 0 0 VSS
port 1 nsew
flabel locali -4520 880 -4270 1040 0 FreeSans 400 0 0 0 I_BIAS
port 6 nsew
flabel locali -5420 -3100 -4990 -2990 0 FreeSans 400 0 0 0 VIN
port 3 nsew
flabel locali -4800 -3100 -4370 -2990 0 FreeSans 400 0 0 0 VIP
port 4 nsew
flabel locali -6070 -3100 -5640 -2990 0 FreeSans 400 0 0 0 VO
port 5 nsew
<< end >>

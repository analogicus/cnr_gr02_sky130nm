magic
tech sky130B
magscale 1 2
timestamp 1713559273
<< metal4 >>
rect -1519 1139 1519 1180
rect -1519 -1139 1263 1139
rect 1499 -1139 1519 1139
rect -1519 -1180 1519 -1139
<< via4 >>
rect 1263 -1139 1499 1139
<< mimcap2 >>
rect -1439 1060 901 1100
rect -1439 -1060 -1399 1060
rect 861 -1060 901 1060
rect -1439 -1100 901 -1060
<< mimcap2contact >>
rect -1399 -1060 861 1060
<< metal5 >>
rect 1221 1139 1541 1181
rect -1423 1060 885 1084
rect -1423 -1060 -1399 1060
rect 861 -1060 885 1060
rect -1423 -1084 885 -1060
rect 1221 -1139 1263 1139
rect 1499 -1139 1541 1139
rect 1221 -1181 1541 -1139
<< properties >>
string FIXED_BBOX -1519 -1180 981 1180
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 11.7 l 11 val 266.025 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

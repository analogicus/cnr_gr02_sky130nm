*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_GR02_lpe.spi
#else
.include ../../../work/xsch/CNR_GR02.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6 keepopinfo noopiter gminsteps=5

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p


*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD  0  dc 1.8

*-----------------------------------------------------------------
* To test OTA
*-----------------------------------------------------------------
*Rin1	in1	vcm1	100
*Rin2	in2	vcm2	100

*vcm1	vcm1	0	dc	.7
*vcm2	vcm2	0	dc	.7
*vin	in1	in2	sin(0	10m	1K)

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VDD VSS CNR_GR02

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.save all
*.save v(VDD) v(VSS) v(xdut.VO) v(xdut.VBJT1) v(xdut.VBJT2) v(xdut.VBJT3) v(xdut.VRO) v(xdut.VRO0) i(vdd) v(xdut.Vb) v(xdut.Vb1)

#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 100n 20u 0

tran 1n 1u 1n

ifdef DEBUG
tran 10p 1n 1p
*quit
#else
dc TEMP -40 125 10
write
quit
#endif

.endc

.end

magic
tech sky130B
magscale 1 2
timestamp 1713555387
<< locali >>
rect 247 4235 17012 4425
rect 16822 3204 17012 4235
rect 4685 3111 5279 3201
rect 4685 3095 5393 3111
rect 5173 3005 5393 3095
rect 12335 2871 12441 2877
rect 10931 2667 10997 2863
rect 11513 2669 11579 2855
rect 12335 2777 12341 2871
rect 12435 2777 12441 2871
rect 10931 2601 11392 2667
rect 11513 2603 12118 2669
rect 11326 1890 11392 2601
rect 12052 1888 12118 2603
rect 12335 2187 12441 2777
rect 12335 2081 12619 2187
rect 12513 2057 12619 2081
rect 12513 1951 12935 2057
rect 11006 1696 11112 1838
rect 11672 1730 11778 1872
rect 11320 1512 11416 1658
rect 11649 1512 11683 1633
rect 11752 1512 11786 1632
rect 12042 1512 12148 1666
rect 12304 1512 12338 1632
rect 11091 1258 12677 1512
rect 12423 152 12677 1258
rect 12422 -40 12946 152
<< viali >>
rect 5393 3005 5499 3111
rect 12341 2777 12435 2871
<< metal1 >>
rect 8428 4236 12676 4340
rect 5387 3111 5505 3123
rect 5387 3005 5393 3111
rect 5499 3005 5603 3111
rect 5709 3005 5715 3111
rect 12335 3045 12441 3051
rect 5387 2993 5505 3005
rect 12335 2871 12441 2939
rect 12335 2777 12341 2871
rect 12435 2777 12441 2871
rect 12335 2765 12441 2777
rect 12572 2592 12676 4236
rect 12572 2488 12926 2592
rect 11570 1750 11872 1800
<< via1 >>
rect 5603 3005 5709 3111
rect 12335 2939 12441 3045
<< metal2 >>
rect 5603 3111 5709 3117
rect 5709 3045 9645 3111
rect 5709 3005 12335 3045
rect 5603 2999 5709 3005
rect 9539 2939 12335 3005
rect 12441 2939 12447 3045
use COMP  COMP_0 
timestamp 1713519326
transform 0 1 15962 -1 0 -2716
box -6200 -3190 -2588 1050
use M6  M6_0 
timestamp 1713519460
transform 0 1 11390 -1 0 1777
box -276 -329 276 329
use M6  M6_1
timestamp 1713519460
transform 0 -1 12045 -1 0 1776
box -276 -329 276 329
use P16  P16_0
timestamp 1713551957
transform 1 0 0 0 1 0
box 0 0 12400 4344
<< end >>

*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/RPLY_EX0_lpe.spi
#else
.include ../../../work/xsch/RPLY_EX0.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TEMP=40 GMIN=1e-15 reltol=1e-6 abstol=1e-6 keepopinfo noopiter gminsteps=5

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD  0  dc 1.8
Vrst rst 0 pwl 0 1.8 10u 1.8 10.01u 0

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VDD VSS rst RPLY_EX0

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.save v(VDD) v(VSS) v(xdut.VO) v(xdut.VBJT1) v(xdut.VBJT2) v(xdut.VBJT3) v(xdut.VRO) v(xdut.VRO0) i(vdd) v(xdut.Vb) v(xdut.Vb1) v(xdut.Vn1) v(xdut.Vn2) v(rst) v(xdut.Vop) v(xdut.Vn20) v(dt)

#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
set file = "tdiff.txt"
unset askquit

optran 0 0 0 100n 20u 0

foreach vtemp -40 -30 -20 -10 0 10 20 30 40 50 60 70 80 90 100 110 120
  option temp=$vtemp
  tran 100n 300u
  meas tran tdiff_$vtemp TRIG V(rst) VAL=0.5 FALL=1 TARG V(xdut.Vop) VAL=.5 FALL=1 >> $file
  write {cicname}_$vtemp
end

let vro0= v(xdut.vro0)
let vref=v(xdut.VRO0)-v(xdut.VBJT2)
let vd= v(xdut.VBJT1)-v(xdut.VRO0)
let W_vdd=i(vdd)*1.8 
let vo=v(xdut.VO)
let vb=v(xdut.Vb)

write
quit
#endif

.endc

.end

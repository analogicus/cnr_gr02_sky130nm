** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/OP_AMP_TESTER_SKY130NM/OP_AMP_TESTER.sch
**.subckt OP_AMP_TESTER VSS VDD_1V8 VIN VIP
*.ipin VSS
*.ipin VDD_1V8
*.ipin VIN
*.ipin VIP
x1 net2 net3 VSS VSS CNRATR_NCH_4C2F0
x2 net3 net3 VSS VSS CNRATR_NCH_4C2F0
x3 net2 VIN net1 net1 CNRATR_PCH_4C4F0
x4 net3 VIP net1 net1 CNRATR_PCH_4C4F0
x5 net1 net5 VDD_1V8 VDD_1V8 CNRATR_PCH_4C4F0
x6 net4 net5 VDD_1V8 net7 CNRATR_PCH_4C4F0
x7 net4 net3 VSS net8 CNRATR_NCH_4C2F0
x8 net6 net5 VDD_1V8 VDD_1V8 CNRATR_PCH_4C4F0
R1 net6 VSS 1k m=1
V1 net4 VSS 0
**** begin user architecture code



* ngspice commands
.include corner.spi



**** end user architecture code
**.ends

* expanding   symbol:  CNR_ATR_SKY130NM/CNRATR_NCH_4C2F0.sym # of pins=4
** sym_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_4C2F0.sym
** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_4C2F0.sch
.subckt CNRATR_NCH_4C2F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.54 W=3.84 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  CNR_ATR_SKY130NM/CNRATR_PCH_4C4F0.sym # of pins=4
** sym_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_4C4F0.sym
** sch_path: /home/solheim22/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_4C4F0.sch
.subckt CNRATR_PCH_4C4F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=1.26 W=3.84 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end

magic
tech sky130B
magscale 1 2
timestamp 1713176887
<< checkpaint >>
rect 7214 5184 16723 5185
rect 7214 5183 23443 5184
rect 7214 5182 30163 5183
rect 7214 5181 36883 5182
rect 7214 5180 43603 5181
rect 7214 5178 50323 5180
rect 7214 -38 59494 5178
rect 6364 -3496 59494 -38
rect 7214 -3497 59494 -3496
rect 13934 -3498 59494 -3497
rect 20654 -3499 59494 -3498
rect 27374 -3500 59494 -3499
rect 34094 -3501 59494 -3500
rect 40814 -3502 59494 -3501
rect 47534 -3503 59494 -3502
rect 50254 -3504 59494 -3503
<< error_s >>
rect 10382 1941 10454 1947
rect 10520 1941 10592 1947
rect 7807 626 7809 1914
rect 10382 1907 10394 1941
rect 10520 1907 10532 1941
rect 10382 1901 10454 1907
rect 10520 1901 10592 1907
rect 10691 1628 10792 1882
rect 9050 1385 9095 1403
rect 9050 1349 9222 1385
rect 9068 753 9222 1349
rect 9607 1315 9642 1349
rect 9608 1296 9642 1315
rect 9268 1247 9340 1253
rect 9406 1247 9478 1253
rect 9268 1213 9280 1247
rect 9406 1213 9418 1247
rect 9268 1207 9340 1213
rect 9406 1207 9478 1213
rect 9068 626 9138 753
rect 9268 719 9340 725
rect 9406 719 9478 725
rect 9268 685 9280 719
rect 9406 685 9418 719
rect 9268 679 9340 685
rect 9406 679 9478 685
rect 9068 600 9129 626
rect 9104 592 9129 600
rect 9627 583 9642 1296
rect 9661 1262 9696 1296
rect 9661 583 9695 1262
rect 9825 1194 9897 1200
rect 9963 1194 10035 1200
rect 9825 1160 9837 1194
rect 9963 1160 9975 1194
rect 9825 1154 9897 1160
rect 9963 1154 10035 1160
rect 9825 666 9897 672
rect 9963 666 10035 672
rect 9825 632 9837 666
rect 9963 632 9975 666
rect 9825 626 9897 632
rect 9963 626 10035 632
rect 9661 549 9676 583
rect 10184 530 10199 1296
rect 10218 530 10252 1350
rect 10382 613 10454 619
rect 10520 613 10592 619
rect 10382 579 10394 613
rect 10520 579 10532 613
rect 10945 594 11046 1628
rect 12079 594 12233 1882
rect 15659 1037 15693 1091
rect 10382 573 10454 579
rect 10520 573 10592 579
rect 10218 496 10233 530
rect 12079 467 12149 594
rect 12079 441 12140 467
rect 12115 433 12140 441
rect 15678 424 15693 1037
rect 15712 1003 15747 1037
rect 15712 424 15746 1003
rect 15873 935 15931 941
rect 15991 935 16049 941
rect 15873 901 15885 935
rect 15991 901 16003 935
rect 15873 895 15931 901
rect 15991 895 16049 901
rect 15873 507 15931 513
rect 15991 507 16049 513
rect 15873 473 15885 507
rect 15991 473 16003 507
rect 15873 467 15931 473
rect 15991 467 16049 473
rect 15712 390 15727 424
rect 16195 371 16210 1037
rect 16229 371 16263 1088
rect 16390 1082 16448 1088
rect 16508 1082 16566 1088
rect 16390 1048 16402 1082
rect 16508 1048 16520 1082
rect 16390 1042 16448 1048
rect 16508 1042 16566 1048
rect 16693 831 16727 885
rect 16390 454 16448 460
rect 16508 454 16566 460
rect 16390 420 16402 454
rect 16508 420 16520 454
rect 16390 414 16448 420
rect 16508 414 16566 420
rect 16229 337 16244 371
rect 16712 318 16727 831
rect 16746 797 16781 831
rect 17289 797 17324 831
rect 16746 318 16780 797
rect 17290 778 17324 797
rect 16746 284 16761 318
rect 17309 265 17324 778
rect 17343 744 17378 778
rect 17343 265 17377 744
rect 17887 693 17921 711
rect 17887 657 17957 693
rect 17904 623 17975 657
rect 18603 623 18638 657
rect 17343 231 17358 265
rect 17904 212 17974 623
rect 18604 604 18638 623
rect 17904 176 17957 212
rect 18623 159 18638 604
rect 18657 570 18692 604
rect 18657 159 18691 570
rect 18657 125 18672 159
rect 2084 -944 2119 -910
rect 2587 -944 2622 -910
rect 1691 -1059 1763 -1053
rect 1829 -1059 1901 -1053
rect 1527 -1086 1561 -1068
rect 26 -1156 1412 -1122
rect -51 -1636 -36 -1156
rect -17 -1183 18 -1156
rect 79 -1177 665 -1156
rect 79 -1183 761 -1177
rect -17 -1583 17 -1183
rect 66 -1200 200 -1190
rect 94 -1224 228 -1218
rect 727 -1224 761 -1183
rect 94 -1228 674 -1224
rect 106 -1258 674 -1228
rect 159 -1285 327 -1258
rect 417 -1285 585 -1258
rect 44 -1296 51 -1292
rect 63 -1296 78 -1292
rect 727 -1296 744 -1245
rect 748 -1296 761 -1224
rect 32 -1400 84 -1296
rect 97 -1323 112 -1319
rect 91 -1324 112 -1323
rect 90 -1335 131 -1324
rect 344 -1335 389 -1324
rect 602 -1335 647 -1324
rect 91 -1400 131 -1335
rect 32 -1481 78 -1400
rect 97 -1431 131 -1400
rect 355 -1431 389 -1335
rect 613 -1431 647 -1335
rect 97 -1447 112 -1431
rect 327 -1481 365 -1443
rect 585 -1481 623 -1443
rect 32 -1496 71 -1481
rect 159 -1496 365 -1481
rect 417 -1496 623 -1481
rect 44 -1500 51 -1496
rect 159 -1500 327 -1496
rect 417 -1500 585 -1496
rect 143 -1515 343 -1500
rect 401 -1515 601 -1500
rect 200 -1521 339 -1515
rect 405 -1521 597 -1515
rect 200 -1534 367 -1528
rect 377 -1534 625 -1528
rect 727 -1534 761 -1296
rect 109 -1549 635 -1534
rect 90 -1568 690 -1549
rect 748 -1582 761 -1534
rect 727 -1583 761 -1582
rect -17 -1617 761 -1583
rect -51 -1651 795 -1636
rect 1491 -1670 1561 -1086
rect 1691 -1093 1703 -1059
rect 1829 -1093 1841 -1059
rect 1691 -1099 1763 -1093
rect 1829 -1099 1901 -1093
rect 1691 -1587 1763 -1581
rect 1829 -1587 1901 -1581
rect 1691 -1621 1703 -1587
rect 1829 -1621 1841 -1587
rect 1691 -1627 1763 -1621
rect 1829 -1627 1901 -1621
rect 1491 -1706 1544 -1670
rect 2050 -1723 2065 -957
rect 2084 -1723 2118 -944
rect 2588 -963 2622 -944
rect 2248 -1012 2320 -1006
rect 2386 -1012 2458 -1006
rect 2248 -1046 2260 -1012
rect 2386 -1046 2398 -1012
rect 2248 -1052 2320 -1046
rect 2386 -1052 2458 -1046
rect 2248 -1640 2320 -1634
rect 2386 -1640 2458 -1634
rect 2248 -1674 2260 -1640
rect 2386 -1674 2398 -1640
rect 2248 -1680 2320 -1674
rect 2386 -1680 2458 -1674
rect 2084 -1757 2099 -1723
rect 2607 -1776 2622 -963
rect 2641 -997 2676 -963
rect 3144 -997 3179 -963
rect 2641 -1776 2675 -997
rect 3145 -1016 3179 -997
rect 2805 -1065 2877 -1059
rect 2943 -1065 3015 -1059
rect 2805 -1099 2817 -1065
rect 2943 -1099 2955 -1065
rect 2805 -1105 2877 -1099
rect 2943 -1105 3015 -1099
rect 2805 -1693 2877 -1687
rect 2943 -1693 3015 -1687
rect 2805 -1727 2817 -1693
rect 2943 -1727 2955 -1693
rect 2805 -1733 2877 -1727
rect 2943 -1733 3015 -1727
rect 2641 -1810 2656 -1776
rect 3164 -1829 3179 -1016
rect 3198 -1050 3233 -1016
rect 3198 -1829 3232 -1050
rect 3362 -1118 3434 -1112
rect 3500 -1118 3572 -1112
rect 3362 -1152 3374 -1118
rect 3500 -1152 3512 -1118
rect 3362 -1158 3434 -1152
rect 3500 -1158 3572 -1152
rect 7103 -1315 7138 -1281
rect 6546 -1357 6581 -1339
rect 6510 -1362 6581 -1357
rect 3702 -1469 3736 -1415
rect 5749 -1427 5784 -1416
rect 4516 -1469 4569 -1434
rect 3362 -1746 3434 -1740
rect 3500 -1746 3572 -1740
rect 3362 -1780 3374 -1746
rect 3500 -1780 3512 -1746
rect 3362 -1786 3434 -1780
rect 3500 -1786 3572 -1780
rect 3198 -1863 3213 -1829
rect 3721 -1882 3736 -1469
rect 3755 -1503 3790 -1469
rect 4498 -1470 4569 -1469
rect 3755 -1882 3789 -1503
rect 4516 -1504 4587 -1470
rect 3755 -1916 3770 -1882
rect 4516 -1935 4586 -1504
rect 4516 -1971 4569 -1935
rect 5715 -1988 5730 -1470
rect 5749 -1988 5783 -1427
rect 5749 -2022 5764 -1988
rect 6510 -2041 6580 -1362
rect 6710 -1430 6782 -1424
rect 6848 -1430 6920 -1424
rect 6710 -1464 6722 -1430
rect 6848 -1464 6860 -1430
rect 6710 -1470 6782 -1464
rect 6848 -1470 6920 -1464
rect 6710 -1958 6782 -1952
rect 6848 -1958 6920 -1952
rect 6710 -1992 6722 -1958
rect 6848 -1992 6860 -1958
rect 6710 -1998 6782 -1992
rect 6848 -1998 6920 -1992
rect 6510 -2077 6563 -2041
rect 7069 -2094 7084 -1328
rect 7103 -2094 7137 -1315
rect 7267 -1383 7339 -1377
rect 7405 -1383 7477 -1377
rect 7267 -1417 7279 -1383
rect 7405 -1417 7417 -1383
rect 7267 -1423 7339 -1417
rect 7405 -1423 7477 -1417
rect 7267 -2011 7339 -2005
rect 7405 -2011 7477 -2005
rect 7267 -2045 7279 -2011
rect 7405 -2045 7417 -2011
rect 7267 -2051 7339 -2045
rect 7405 -2051 7477 -2045
rect 7103 -2128 7118 -2094
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
use COMP  x2
timestamp 0
transform 1 0 0 0 1 600
box 0 0 1 1
use sky130_fd_pr__cap_mim_m3_2_3HBNLG  XC1
timestamp 0
transform 1 0 11823 0 1 844
box -3349 -3081 3371 3081
use sky130_fd_pr__cap_mim_m3_2_3HBNLG  XC2
timestamp 0
transform 1 0 18543 0 1 843
box -3349 -3081 3371 3081
use sky130_fd_pr__cap_mim_m3_2_3HBNLG  XC3
timestamp 0
transform 1 0 25263 0 1 842
box -3349 -3081 3371 3081
use sky130_fd_pr__cap_mim_m3_2_3HBNLG  XC4
timestamp 0
transform 1 0 31983 0 1 841
box -3349 -3081 3371 3081
use sky130_fd_pr__cap_mim_m3_2_3HBNLG  XC5
timestamp 0
transform 1 0 38703 0 1 840
box -3349 -3081 3371 3081
use sky130_fd_pr__cap_mim_m3_2_3HBNLG  XC6
timestamp 0
transform 1 0 45423 0 1 839
box -3349 -3081 3371 3081
use sky130_fd_pr__cap_mim_m3_2_4PHTN9  XC7
timestamp 0
transform 1 0 50143 0 1 -1162
box -1349 -1081 1371 1081
use sky130_fd_pr__cap_mim_m3_2_3HBNLG  XC8
timestamp 0
transform 1 0 54863 0 1 837
box -3349 -3081 3371 3081
use sky130_fd_pr__pfet_01v8_JMC8WZ  XM1
timestamp 0
transform 1 0 15961 0 1 704
box -285 -369 285 369
use sky130_fd_pr__pfet_01v8_JMP7WZ  XM2
timestamp 0
transform 1 0 16478 0 1 751
box -285 -469 285 469
use sky130_fd_pr__pfet_01v8_XPC8Y6  XM3
timestamp 0
transform 1 0 17035 0 1 548
box -325 -319 325 319
use sky130_fd_pr__pfet_01v8_XPC8Y6  XM4
timestamp 0
transform 1 0 17632 0 1 495
box -325 -319 325 319
use sky130_fd_pr__nfet_01v8_U7AL37  XM5
timestamp 0
transform 1 0 18289 0 1 408
box -385 -285 385 285
use sky130_fd_pr__nfet_01v8_U7AL37  XM6
timestamp 0
transform 1 0 19006 0 1 355
box -385 -285 385 285
use sky130_fd_pr__nfet_01v8_ZYANF2  XM7
timestamp 0
transform 1 0 372 0 1 -1383
box -425 -270 425 270
use sky130_fd_pr__nfet_01v8_RFVHWA  XM8
timestamp 0
transform 1 0 719 0 1 -1396
box -825 -310 825 310
use sky130_fd_pr__pfet_01v8_XPP79A  XM9
timestamp 0
transform 1 0 1796 0 1 -1340
box -305 -419 305 419
use sky130_fd_pr__pfet_01v8_TMP79A  XM10
timestamp 0
transform 1 0 2353 0 1 -1343
box -305 -469 305 469
use sky130_fd_pr__pfet_01v8_TMP79A  XM11
timestamp 0
transform 1 0 2910 0 1 -1396
box -305 -469 305 469
use sky130_fd_pr__pfet_01v8_XPP79A  XM12
timestamp 0
transform 1 0 9373 0 1 966
box -305 -419 305 419
use sky130_fd_pr__pfet_01v8_XPP79A  XM13
timestamp 0
transform 1 0 9930 0 1 913
box -305 -419 305 419
use sky130_fd_pr__pfet_01v8_XPB89A  XM14
timestamp 0
transform 1 0 10487 0 1 1260
box -305 -819 305 819
use sky130_fd_pr__pfet_01v8_XPP79A  XM15
timestamp 0
transform 1 0 6815 0 1 -1711
box -305 -419 305 419
use sky130_fd_pr__pfet_01v8_CQBZVD  XM16
timestamp 0
transform 1 0 13904 0 1 1357
box -1825 -969 1825 969
use sky130_fd_pr__pfet_01v8_TMP79A  XM17
timestamp 0
transform 1 0 3467 0 1 -1449
box -305 -469 305 469
use sky130_fd_pr__pfet_01v8_TMP79A  XM18
timestamp 0
transform 1 0 7372 0 1 -1714
box -305 -469 305 469
use sky130_fd_pr__pfet_01v8_FQU9VM  XM19
timestamp 0
transform 1 0 8049 0 1 -1767
box -425 -469 425 469
use sky130_fd_pr__pfet_01v8_FQE7VM  XM21
timestamp 0
transform 1 0 4144 0 1 -1702
box -425 -269 425 269
use sky130_fd_pr__nfet_01v8_UTAWZB  XM22
timestamp 0
transform 1 0 5141 0 1 -1729
box -625 -295 625 295
use sky130_fd_pr__nfet_01v8_QGMQ49  XM27
timestamp 0
transform 1 0 6138 0 1 -1717
box -425 -360 425 360
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ1 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1705202102
transform 1 0 7781 0 1 600
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ2
array 0 5 1288 0 0 1288
timestamp 1705202102
transform 1 0 1 0 1 600
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ3
timestamp 1705202102
transform 1 0 10792 0 1 441
box 0 0 1340 1340
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD_1V8
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 rst
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 LPO
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 LPI
port 4 nsew
<< end >>

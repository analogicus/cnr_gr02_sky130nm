magic
tech sky130B
magscale 1 2
timestamp 1713546649
<< nwell >>
rect 3960 3042 6445 4120
<< locali >>
rect 5946 4129 6214 4130
rect 4902 4085 6214 4129
rect 4902 4084 5991 4085
rect 4902 4022 4947 4084
rect 5417 4030 5462 4084
rect 5946 4020 5991 4084
rect 4721 3872 4819 3906
rect 4597 3613 4631 3727
rect 4721 3679 4755 3872
rect 4878 3679 4923 3748
rect 5459 3679 5504 3754
rect 5878 3679 5923 3752
rect 6169 3679 6214 4085
rect 6297 4062 6331 4221
rect 3546 2141 3660 3206
rect 4685 3095 4791 3679
rect 4878 3634 6214 3679
rect 6297 3559 6331 3716
rect 5864 3525 6331 3559
rect 5864 3446 5898 3525
rect 3874 2420 4306 2576
rect 5176 2568 5608 2724
rect 5176 2246 5608 2402
rect 3876 2064 4308 2220
rect 4050 1796 5194 1912
rect 5864 1635 5898 1718
rect 6487 1635 6521 1753
rect 7185 1635 7219 1753
rect 7971 1635 8005 1755
rect 8753 1635 8787 1755
rect 9126 1635 9160 1718
rect 5864 1601 9160 1635
rect 7500 1258 10405 1512
<< viali >>
rect 4685 2989 4791 3095
rect 3546 2027 3660 2141
<< metal1 >>
rect 4310 3682 4362 3928
rect 6046 3866 6252 3918
rect 3015 3630 4362 3682
rect 5961 3588 6007 3589
rect 6200 3588 6252 3866
rect 5961 3536 6252 3588
rect 5961 3366 6007 3536
rect 4483 3041 4537 3252
rect 3093 2987 4537 3041
rect 4673 3095 4803 3101
rect 4673 2989 4685 3095
rect 4791 2989 4803 3095
rect 4673 2983 4803 2989
rect 4685 2813 4791 2983
rect 3877 2707 4791 2813
rect 3534 2141 3672 2147
rect 3534 2027 3546 2141
rect 3660 2027 3672 2141
rect 5176 2036 5827 2106
rect 3534 2021 3672 2027
rect 3546 1615 3660 2021
rect 5246 803 5360 1674
rect 5757 1518 5827 2036
rect 5757 1447 8359 1518
rect 8288 781 8359 1447
use M14  M14_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713520534
transform 0 1 5443 -1 0 3889
box -305 -919 305 1002
use M16  M16_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713520667
transform 0 -1 7512 -1 0 2582
box -996 -1684 996 1684
use M27  M27_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713522689
transform 0 1 11689 -1 0 3222
box -296 -479 296 479
use p7  p7_0
timestamp 1713528272
transform 1 0 12 0 1 1416
box -12 -1416 7768 2830
use Q2  Q2_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713441746
transform 1 0 2 0 1 -600
box 7780 600 9120 1940
use sky130_fd_pr__res_high_po_0p35_CMWQMJ  sky130_fd_pr__res_high_po_0p35_CMWQMJ_0
timestamp 0
transform 0 1 4742 -1 0 2403
box -533 -1032 533 1032
use sky130_fd_pr__res_high_po_0p35_N7UQCW  sky130_fd_pr__res_high_po_0p35_N7UQCW_0
timestamp 0
transform 0 1 4449 -1 0 1649
box -201 -1237 201 1237
<< end >>

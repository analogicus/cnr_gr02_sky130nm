magic
tech sky130B
magscale 1 2
timestamp 1713542901
<< locali >>
rect 5946 4129 6214 4130
rect 4902 4085 6214 4129
rect 4902 4084 5991 4085
rect 4902 4022 4947 4084
rect 5417 4030 5462 4084
rect 5946 4020 5991 4084
rect 4597 3613 4631 3727
rect 4878 3679 4923 3748
rect 5459 3679 5504 3754
rect 5878 3679 5923 3752
rect 6169 3679 6214 4085
rect 6297 4062 6331 4221
rect 4878 3634 6214 3679
rect 3546 2141 3660 3206
<< viali >>
rect 3546 2027 3660 2141
<< metal1 >>
rect 4310 3682 4362 3928
rect 3015 3630 4362 3682
rect 4483 3041 4537 3252
rect 3093 2987 4537 3041
rect 3534 2141 3672 2147
rect 3534 2027 3546 2141
rect 3660 2027 3672 2141
rect 3534 2021 3672 2027
rect 3546 1615 3660 2021
rect 5246 803 5360 1674
use M14  M14_0 ~/lpro/temp_to_current_temp1_layout1/rply_ex0_sky130nm/design/RPLY_EX0_SKY130NM/mag
timestamp 1713520534
transform 0 1 5443 -1 0 3889
box -305 -919 305 1002
use p7  p7_0
timestamp 1713528272
transform 1 0 12 0 1 1416
box -12 -1416 7768 2830
use sky130_fd_pr__res_high_po_0p35_N7UQCW  sky130_fd_pr__res_high_po_0p35_N7UQCW_0
timestamp 0
transform 0 1 4449 -1 0 1649
box -201 -1237 201 1237
<< end >>

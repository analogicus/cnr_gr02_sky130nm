magic
tech sky130B
magscale 1 2
timestamp 1713258222
<< error_p >>
rect -105 681 -33 687
rect 33 681 105 687
rect -105 647 -93 681
rect 33 647 45 681
rect -105 641 -33 647
rect 33 641 105 647
rect -105 -647 -33 -641
rect 33 -647 105 -641
rect -105 -681 -93 -647
rect 33 -681 45 -647
rect -105 -687 -33 -681
rect 33 -687 105 -681
<< nwell >>
rect -305 -819 305 819
<< pmos >>
rect -109 -600 -29 600
rect 29 -600 109 600
<< pdiff >>
rect -167 588 -109 600
rect -167 -588 -155 588
rect -121 -588 -109 588
rect -167 -600 -109 -588
rect -29 588 29 600
rect -29 -588 -17 588
rect 17 -588 29 588
rect -29 -600 29 -588
rect 109 588 167 600
rect 109 -588 121 588
rect 155 -588 167 588
rect 109 -600 167 -588
<< pdiffc >>
rect -155 -588 -121 588
rect -17 -588 17 588
rect 121 -588 155 588
<< nsubdiff >>
rect -269 749 -173 783
rect 173 749 269 783
rect -269 687 -235 749
rect 235 687 269 749
rect -269 -749 -235 -687
rect 235 -749 269 -687
rect -269 -783 -173 -749
rect 173 -783 269 -749
<< nsubdiffcont >>
rect -173 749 173 783
rect -269 -687 -235 687
rect 235 -687 269 687
rect -173 -783 173 -749
<< poly >>
rect -109 681 -29 697
rect -109 647 -93 681
rect -45 647 -29 681
rect -109 600 -29 647
rect 29 681 109 697
rect 29 647 45 681
rect 93 647 109 681
rect 29 600 109 647
rect -109 -647 -29 -600
rect -109 -681 -93 -647
rect -45 -681 -29 -647
rect -109 -697 -29 -681
rect 29 -647 109 -600
rect 29 -681 45 -647
rect 93 -681 109 -647
rect 29 -697 109 -681
<< polycont >>
rect -93 647 -45 681
rect 45 647 93 681
rect -93 -681 -45 -647
rect 45 -681 93 -647
<< locali >>
rect -269 749 -173 783
rect 173 749 269 783
rect -269 687 -235 749
rect 235 687 269 749
rect -109 647 -93 681
rect -45 647 -29 681
rect 29 647 45 681
rect 93 647 109 681
rect -155 588 -121 604
rect -155 -604 -121 -588
rect -17 588 17 604
rect -17 -604 17 -588
rect 121 588 155 604
rect 121 -604 155 -588
rect -109 -681 -93 -647
rect -45 -681 -29 -647
rect 29 -681 45 -647
rect 93 -681 109 -647
rect -269 -749 -235 -687
rect 235 -749 269 -687
rect -269 -783 -173 -749
rect 173 -783 269 -749
<< viali >>
rect -93 647 -45 681
rect 45 647 93 681
rect -155 -588 -121 588
rect -17 -588 17 588
rect 121 -588 155 588
rect -93 -681 -45 -647
rect 45 -681 93 -647
<< metal1 >>
rect -105 681 -33 687
rect -105 647 -93 681
rect -45 647 -33 681
rect -105 641 -33 647
rect 33 681 105 687
rect 33 647 45 681
rect 93 647 105 681
rect 33 641 105 647
rect -161 588 -115 600
rect -161 -588 -155 588
rect -121 -588 -115 588
rect -161 -600 -115 -588
rect -23 588 23 600
rect -23 -588 -17 588
rect 17 -588 23 588
rect -23 -600 23 -588
rect 115 588 161 600
rect 115 -588 121 588
rect 155 -588 161 588
rect 115 -600 161 -588
rect -105 -647 -33 -641
rect -105 -681 -93 -647
rect -45 -681 -33 -647
rect -105 -687 -33 -681
rect 33 -647 105 -641
rect 33 -681 45 -647
rect 93 -681 105 -647
rect 33 -687 105 -681
<< properties >>
string FIXED_BBOX -252 -766 252 766
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.0 l 0.4 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130B
magscale 1 2
timestamp 1713553862
<< locali >>
rect 10931 2667 10997 2863
rect 11513 2669 11579 2855
rect 10931 2601 11392 2667
rect 11513 2603 12118 2669
rect 11326 1890 11392 2601
rect 12052 1888 12118 2603
rect 11006 1696 11112 1838
rect 11672 1730 11778 1872
rect 11320 1512 11416 1658
rect 11649 1512 11683 1633
rect 11752 1512 11786 1632
rect 12042 1512 12148 1666
rect 12304 1512 12338 1632
rect 11091 1258 12677 1512
<< metal1 >>
rect 11570 1750 11872 1800
use M6  M6_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713519460
transform 0 1 11390 -1 0 1777
box -276 -329 276 329
use M6  M6_1
timestamp 1713519460
transform 0 -1 12045 -1 0 1776
box -276 -329 276 329
use P16  P16_0
timestamp 1713551957
transform 1 0 0 0 1 0
box 0 0 12400 4344
<< end >>

magic
tech sky130B
magscale 1 2
timestamp 1713518682
<< pwell >>
rect -396 -349 396 349
<< nmos >>
rect -200 -201 200 139
<< ndiff >>
rect -258 127 -200 139
rect -258 -189 -246 127
rect -212 -189 -200 127
rect -258 -201 -200 -189
rect 200 127 258 139
rect 200 -189 212 127
rect 246 -189 258 127
rect 200 -201 258 -189
<< ndiffc >>
rect -246 -189 -212 127
rect 212 -189 246 127
<< psubdiff >>
rect -326 279 -264 313
rect 264 279 326 313
rect -326 -313 -264 -279
rect 264 -313 326 -279
<< psubdiffcont >>
rect -264 279 264 313
rect -264 -313 264 -279
<< poly >>
rect -373 -228 -317 228
rect -200 211 200 227
rect -200 177 -184 211
rect 184 177 200 211
rect -200 139 200 177
rect -200 -227 200 -201
rect 323 -226 379 230
<< polycont >>
rect -184 177 184 211
<< locali >>
rect -280 279 -264 313
rect 264 279 280 313
rect -200 177 -184 211
rect 184 177 200 211
rect -246 127 -212 143
rect -246 -205 -212 -189
rect 212 127 246 143
rect 212 -205 246 -189
rect -280 -313 -264 -279
rect 264 -313 280 -279
<< viali >>
rect -184 177 184 211
rect -246 -189 -212 127
rect 212 -189 246 127
<< metal1 >>
rect -196 211 196 217
rect -196 177 -184 211
rect 184 177 196 211
rect -196 171 196 177
rect -252 127 -206 139
rect -252 -189 -246 127
rect -212 -189 -206 127
rect -252 -201 -206 -189
rect 206 127 252 139
rect 206 -189 212 127
rect 246 -189 252 127
rect 206 -201 252 -189
<< properties >>
string FIXED_BBOX -343 -296 343 296
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.7 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

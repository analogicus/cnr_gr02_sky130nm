magic
tech sky130B
magscale 1 2
timestamp 1713527212
<< nwell >>
rect 806 1626 3268 2698
<< locali >>
rect 1915 2784 3429 2830
rect 2052 2572 2086 2784
rect 2527 2529 2573 2784
rect 3114 2572 3148 2784
rect 1924 2426 2062 2504
rect 2512 1934 2606 2390
rect 3114 2179 3148 2364
rect 3114 2145 3223 2179
rect 3189 1963 3223 2145
rect 1822 1834 1960 1912
rect 1734 0 3870 96
<< viali >>
rect 641 1577 683 1619
<< metal1 >>
rect 3003 2266 3055 2444
rect 1814 2214 3055 2266
rect 3081 1625 3135 1840
rect 629 1619 3135 1625
rect 629 1577 641 1619
rect 683 1577 3135 1619
rect 629 1571 3135 1577
use M9  M9_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713524830
transform 0 1 2600 -1 0 2468
box -236 -584 236 584
use M10  M10_0 ~/aicex/ip/cnr_gr02_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1713518505
transform 0 1 2580 -1 0 1864
box -236 -684 236 684
use p4  p4_0
timestamp 1713525798
transform 1 0 0 0 1 0
box 0 0 1980 2830
<< end >>

*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/COMP_lpe.spi
#else
.include ../../../work/xsch/COMP.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD  0  dc 1.8
I_BIAS 0 I_TEST dc 5u
VIP VIP 0 dc 0.9
VIN VIN 0 SIN(0.9 0.9 10 0 0)
VNY I_TEST I_BIAS dc 0
*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VSS VDD VIN VIP VO I_BIAS COMP

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 10n 10u 0
tran 100u 300m 1n
write
quit


.endc

.end
